`timescale 1ns/10ps
module controller(
	clk,
	rst,
	all_layer_set_done,
);