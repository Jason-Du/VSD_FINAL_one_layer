# 
#              Synchronous Dual Port SRAM Compiler 
# 
#                    UMC 0.18um Generic Logic Process 
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : word64
#       Words            : 64
#       Bits             : 16
#       Byte-Write       : 8
#       Aspect Ratio     : 1
#       Output Loading   : 0.5  (pf)
#       Data Slew        : 0.5  (ns)
#       CK Slew          : 0.5  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2021/01/11 17:17:22
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO word64
CLASS BLOCK ;
FOREIGN word64 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 3547.640 BY 179.760 ;
SYMMETRY x y r90 ;
SITE core ;
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal5 ;
  RECT 3546.520 168.340 3547.640 171.580 ;
  LAYER metal4 ;
  RECT 3546.520 168.340 3547.640 171.580 ;
  LAYER metal3 ;
  RECT 3546.520 168.340 3547.640 171.580 ;
  LAYER metal2 ;
  RECT 3546.520 168.340 3547.640 171.580 ;
  LAYER metal1 ;
  RECT 3546.520 168.340 3547.640 171.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3546.520 129.140 3547.640 132.380 ;
  LAYER metal4 ;
  RECT 3546.520 129.140 3547.640 132.380 ;
  LAYER metal3 ;
  RECT 3546.520 129.140 3547.640 132.380 ;
  LAYER metal2 ;
  RECT 3546.520 129.140 3547.640 132.380 ;
  LAYER metal1 ;
  RECT 3546.520 129.140 3547.640 132.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3546.520 121.300 3547.640 124.540 ;
  LAYER metal4 ;
  RECT 3546.520 121.300 3547.640 124.540 ;
  LAYER metal3 ;
  RECT 3546.520 121.300 3547.640 124.540 ;
  LAYER metal2 ;
  RECT 3546.520 121.300 3547.640 124.540 ;
  LAYER metal1 ;
  RECT 3546.520 121.300 3547.640 124.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3546.520 113.460 3547.640 116.700 ;
  LAYER metal4 ;
  RECT 3546.520 113.460 3547.640 116.700 ;
  LAYER metal3 ;
  RECT 3546.520 113.460 3547.640 116.700 ;
  LAYER metal2 ;
  RECT 3546.520 113.460 3547.640 116.700 ;
  LAYER metal1 ;
  RECT 3546.520 113.460 3547.640 116.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3546.520 105.620 3547.640 108.860 ;
  LAYER metal4 ;
  RECT 3546.520 105.620 3547.640 108.860 ;
  LAYER metal3 ;
  RECT 3546.520 105.620 3547.640 108.860 ;
  LAYER metal2 ;
  RECT 3546.520 105.620 3547.640 108.860 ;
  LAYER metal1 ;
  RECT 3546.520 105.620 3547.640 108.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3546.520 97.780 3547.640 101.020 ;
  LAYER metal4 ;
  RECT 3546.520 97.780 3547.640 101.020 ;
  LAYER metal3 ;
  RECT 3546.520 97.780 3547.640 101.020 ;
  LAYER metal2 ;
  RECT 3546.520 97.780 3547.640 101.020 ;
  LAYER metal1 ;
  RECT 3546.520 97.780 3547.640 101.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3546.520 89.940 3547.640 93.180 ;
  LAYER metal4 ;
  RECT 3546.520 89.940 3547.640 93.180 ;
  LAYER metal3 ;
  RECT 3546.520 89.940 3547.640 93.180 ;
  LAYER metal2 ;
  RECT 3546.520 89.940 3547.640 93.180 ;
  LAYER metal1 ;
  RECT 3546.520 89.940 3547.640 93.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3546.520 50.740 3547.640 53.980 ;
  LAYER metal4 ;
  RECT 3546.520 50.740 3547.640 53.980 ;
  LAYER metal3 ;
  RECT 3546.520 50.740 3547.640 53.980 ;
  LAYER metal2 ;
  RECT 3546.520 50.740 3547.640 53.980 ;
  LAYER metal1 ;
  RECT 3546.520 50.740 3547.640 53.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3546.520 42.900 3547.640 46.140 ;
  LAYER metal4 ;
  RECT 3546.520 42.900 3547.640 46.140 ;
  LAYER metal3 ;
  RECT 3546.520 42.900 3547.640 46.140 ;
  LAYER metal2 ;
  RECT 3546.520 42.900 3547.640 46.140 ;
  LAYER metal1 ;
  RECT 3546.520 42.900 3547.640 46.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3546.520 35.060 3547.640 38.300 ;
  LAYER metal4 ;
  RECT 3546.520 35.060 3547.640 38.300 ;
  LAYER metal3 ;
  RECT 3546.520 35.060 3547.640 38.300 ;
  LAYER metal2 ;
  RECT 3546.520 35.060 3547.640 38.300 ;
  LAYER metal1 ;
  RECT 3546.520 35.060 3547.640 38.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3546.520 27.220 3547.640 30.460 ;
  LAYER metal4 ;
  RECT 3546.520 27.220 3547.640 30.460 ;
  LAYER metal3 ;
  RECT 3546.520 27.220 3547.640 30.460 ;
  LAYER metal2 ;
  RECT 3546.520 27.220 3547.640 30.460 ;
  LAYER metal1 ;
  RECT 3546.520 27.220 3547.640 30.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3546.520 19.380 3547.640 22.620 ;
  LAYER metal4 ;
  RECT 3546.520 19.380 3547.640 22.620 ;
  LAYER metal3 ;
  RECT 3546.520 19.380 3547.640 22.620 ;
  LAYER metal2 ;
  RECT 3546.520 19.380 3547.640 22.620 ;
  LAYER metal1 ;
  RECT 3546.520 19.380 3547.640 22.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3546.520 11.540 3547.640 14.780 ;
  LAYER metal4 ;
  RECT 3546.520 11.540 3547.640 14.780 ;
  LAYER metal3 ;
  RECT 3546.520 11.540 3547.640 14.780 ;
  LAYER metal2 ;
  RECT 3546.520 11.540 3547.640 14.780 ;
  LAYER metal1 ;
  RECT 3546.520 11.540 3547.640 14.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER metal4 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER metal3 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER metal2 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER metal1 ;
  RECT 0.000 168.340 1.120 171.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER metal4 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER metal3 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER metal2 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER metal1 ;
  RECT 0.000 129.140 1.120 132.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER metal4 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER metal3 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER metal2 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER metal1 ;
  RECT 0.000 121.300 1.120 124.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER metal4 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER metal3 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER metal2 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER metal1 ;
  RECT 0.000 113.460 1.120 116.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER metal4 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER metal3 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER metal2 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER metal1 ;
  RECT 0.000 105.620 1.120 108.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER metal4 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER metal3 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER metal2 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER metal1 ;
  RECT 0.000 97.780 1.120 101.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER metal4 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER metal3 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER metal2 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER metal1 ;
  RECT 0.000 89.940 1.120 93.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER metal4 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER metal3 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER metal2 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER metal1 ;
  RECT 0.000 50.740 1.120 53.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER metal4 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER metal3 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER metal2 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER metal1 ;
  RECT 0.000 42.900 1.120 46.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER metal4 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER metal3 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER metal2 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER metal1 ;
  RECT 0.000 35.060 1.120 38.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER metal4 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER metal3 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER metal2 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER metal1 ;
  RECT 0.000 27.220 1.120 30.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER metal4 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER metal3 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER metal2 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER metal1 ;
  RECT 0.000 19.380 1.120 22.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER metal4 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER metal3 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER metal2 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER metal1 ;
  RECT 0.000 11.540 1.120 14.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3531.300 178.640 3534.840 179.760 ;
  LAYER metal4 ;
  RECT 3531.300 178.640 3534.840 179.760 ;
  LAYER metal3 ;
  RECT 3531.300 178.640 3534.840 179.760 ;
  LAYER metal2 ;
  RECT 3531.300 178.640 3534.840 179.760 ;
  LAYER metal1 ;
  RECT 3531.300 178.640 3534.840 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3517.660 178.640 3521.200 179.760 ;
  LAYER metal4 ;
  RECT 3517.660 178.640 3521.200 179.760 ;
  LAYER metal3 ;
  RECT 3517.660 178.640 3521.200 179.760 ;
  LAYER metal2 ;
  RECT 3517.660 178.640 3521.200 179.760 ;
  LAYER metal1 ;
  RECT 3517.660 178.640 3521.200 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3450.700 178.640 3454.240 179.760 ;
  LAYER metal4 ;
  RECT 3450.700 178.640 3454.240 179.760 ;
  LAYER metal3 ;
  RECT 3450.700 178.640 3454.240 179.760 ;
  LAYER metal2 ;
  RECT 3450.700 178.640 3454.240 179.760 ;
  LAYER metal1 ;
  RECT 3450.700 178.640 3454.240 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3437.060 178.640 3440.600 179.760 ;
  LAYER metal4 ;
  RECT 3437.060 178.640 3440.600 179.760 ;
  LAYER metal3 ;
  RECT 3437.060 178.640 3440.600 179.760 ;
  LAYER metal2 ;
  RECT 3437.060 178.640 3440.600 179.760 ;
  LAYER metal1 ;
  RECT 3437.060 178.640 3440.600 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3423.420 178.640 3426.960 179.760 ;
  LAYER metal4 ;
  RECT 3423.420 178.640 3426.960 179.760 ;
  LAYER metal3 ;
  RECT 3423.420 178.640 3426.960 179.760 ;
  LAYER metal2 ;
  RECT 3423.420 178.640 3426.960 179.760 ;
  LAYER metal1 ;
  RECT 3423.420 178.640 3426.960 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3410.400 178.640 3413.940 179.760 ;
  LAYER metal4 ;
  RECT 3410.400 178.640 3413.940 179.760 ;
  LAYER metal3 ;
  RECT 3410.400 178.640 3413.940 179.760 ;
  LAYER metal2 ;
  RECT 3410.400 178.640 3413.940 179.760 ;
  LAYER metal1 ;
  RECT 3410.400 178.640 3413.940 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3396.760 178.640 3400.300 179.760 ;
  LAYER metal4 ;
  RECT 3396.760 178.640 3400.300 179.760 ;
  LAYER metal3 ;
  RECT 3396.760 178.640 3400.300 179.760 ;
  LAYER metal2 ;
  RECT 3396.760 178.640 3400.300 179.760 ;
  LAYER metal1 ;
  RECT 3396.760 178.640 3400.300 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3383.120 178.640 3386.660 179.760 ;
  LAYER metal4 ;
  RECT 3383.120 178.640 3386.660 179.760 ;
  LAYER metal3 ;
  RECT 3383.120 178.640 3386.660 179.760 ;
  LAYER metal2 ;
  RECT 3383.120 178.640 3386.660 179.760 ;
  LAYER metal1 ;
  RECT 3383.120 178.640 3386.660 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3316.160 178.640 3319.700 179.760 ;
  LAYER metal4 ;
  RECT 3316.160 178.640 3319.700 179.760 ;
  LAYER metal3 ;
  RECT 3316.160 178.640 3319.700 179.760 ;
  LAYER metal2 ;
  RECT 3316.160 178.640 3319.700 179.760 ;
  LAYER metal1 ;
  RECT 3316.160 178.640 3319.700 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3302.520 178.640 3306.060 179.760 ;
  LAYER metal4 ;
  RECT 3302.520 178.640 3306.060 179.760 ;
  LAYER metal3 ;
  RECT 3302.520 178.640 3306.060 179.760 ;
  LAYER metal2 ;
  RECT 3302.520 178.640 3306.060 179.760 ;
  LAYER metal1 ;
  RECT 3302.520 178.640 3306.060 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3288.880 178.640 3292.420 179.760 ;
  LAYER metal4 ;
  RECT 3288.880 178.640 3292.420 179.760 ;
  LAYER metal3 ;
  RECT 3288.880 178.640 3292.420 179.760 ;
  LAYER metal2 ;
  RECT 3288.880 178.640 3292.420 179.760 ;
  LAYER metal1 ;
  RECT 3288.880 178.640 3292.420 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3275.860 178.640 3279.400 179.760 ;
  LAYER metal4 ;
  RECT 3275.860 178.640 3279.400 179.760 ;
  LAYER metal3 ;
  RECT 3275.860 178.640 3279.400 179.760 ;
  LAYER metal2 ;
  RECT 3275.860 178.640 3279.400 179.760 ;
  LAYER metal1 ;
  RECT 3275.860 178.640 3279.400 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3262.220 178.640 3265.760 179.760 ;
  LAYER metal4 ;
  RECT 3262.220 178.640 3265.760 179.760 ;
  LAYER metal3 ;
  RECT 3262.220 178.640 3265.760 179.760 ;
  LAYER metal2 ;
  RECT 3262.220 178.640 3265.760 179.760 ;
  LAYER metal1 ;
  RECT 3262.220 178.640 3265.760 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3248.580 178.640 3252.120 179.760 ;
  LAYER metal4 ;
  RECT 3248.580 178.640 3252.120 179.760 ;
  LAYER metal3 ;
  RECT 3248.580 178.640 3252.120 179.760 ;
  LAYER metal2 ;
  RECT 3248.580 178.640 3252.120 179.760 ;
  LAYER metal1 ;
  RECT 3248.580 178.640 3252.120 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3181.620 178.640 3185.160 179.760 ;
  LAYER metal4 ;
  RECT 3181.620 178.640 3185.160 179.760 ;
  LAYER metal3 ;
  RECT 3181.620 178.640 3185.160 179.760 ;
  LAYER metal2 ;
  RECT 3181.620 178.640 3185.160 179.760 ;
  LAYER metal1 ;
  RECT 3181.620 178.640 3185.160 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3167.980 178.640 3171.520 179.760 ;
  LAYER metal4 ;
  RECT 3167.980 178.640 3171.520 179.760 ;
  LAYER metal3 ;
  RECT 3167.980 178.640 3171.520 179.760 ;
  LAYER metal2 ;
  RECT 3167.980 178.640 3171.520 179.760 ;
  LAYER metal1 ;
  RECT 3167.980 178.640 3171.520 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3154.960 178.640 3158.500 179.760 ;
  LAYER metal4 ;
  RECT 3154.960 178.640 3158.500 179.760 ;
  LAYER metal3 ;
  RECT 3154.960 178.640 3158.500 179.760 ;
  LAYER metal2 ;
  RECT 3154.960 178.640 3158.500 179.760 ;
  LAYER metal1 ;
  RECT 3154.960 178.640 3158.500 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3141.320 178.640 3144.860 179.760 ;
  LAYER metal4 ;
  RECT 3141.320 178.640 3144.860 179.760 ;
  LAYER metal3 ;
  RECT 3141.320 178.640 3144.860 179.760 ;
  LAYER metal2 ;
  RECT 3141.320 178.640 3144.860 179.760 ;
  LAYER metal1 ;
  RECT 3141.320 178.640 3144.860 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3127.680 178.640 3131.220 179.760 ;
  LAYER metal4 ;
  RECT 3127.680 178.640 3131.220 179.760 ;
  LAYER metal3 ;
  RECT 3127.680 178.640 3131.220 179.760 ;
  LAYER metal2 ;
  RECT 3127.680 178.640 3131.220 179.760 ;
  LAYER metal1 ;
  RECT 3127.680 178.640 3131.220 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3116.520 178.640 3120.060 179.760 ;
  LAYER metal4 ;
  RECT 3116.520 178.640 3120.060 179.760 ;
  LAYER metal3 ;
  RECT 3116.520 178.640 3120.060 179.760 ;
  LAYER metal2 ;
  RECT 3116.520 178.640 3120.060 179.760 ;
  LAYER metal1 ;
  RECT 3116.520 178.640 3120.060 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3047.080 178.640 3050.620 179.760 ;
  LAYER metal4 ;
  RECT 3047.080 178.640 3050.620 179.760 ;
  LAYER metal3 ;
  RECT 3047.080 178.640 3050.620 179.760 ;
  LAYER metal2 ;
  RECT 3047.080 178.640 3050.620 179.760 ;
  LAYER metal1 ;
  RECT 3047.080 178.640 3050.620 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3034.060 178.640 3037.600 179.760 ;
  LAYER metal4 ;
  RECT 3034.060 178.640 3037.600 179.760 ;
  LAYER metal3 ;
  RECT 3034.060 178.640 3037.600 179.760 ;
  LAYER metal2 ;
  RECT 3034.060 178.640 3037.600 179.760 ;
  LAYER metal1 ;
  RECT 3034.060 178.640 3037.600 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3020.420 178.640 3023.960 179.760 ;
  LAYER metal4 ;
  RECT 3020.420 178.640 3023.960 179.760 ;
  LAYER metal3 ;
  RECT 3020.420 178.640 3023.960 179.760 ;
  LAYER metal2 ;
  RECT 3020.420 178.640 3023.960 179.760 ;
  LAYER metal1 ;
  RECT 3020.420 178.640 3023.960 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3006.780 178.640 3010.320 179.760 ;
  LAYER metal4 ;
  RECT 3006.780 178.640 3010.320 179.760 ;
  LAYER metal3 ;
  RECT 3006.780 178.640 3010.320 179.760 ;
  LAYER metal2 ;
  RECT 3006.780 178.640 3010.320 179.760 ;
  LAYER metal1 ;
  RECT 3006.780 178.640 3010.320 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2993.760 178.640 2997.300 179.760 ;
  LAYER metal4 ;
  RECT 2993.760 178.640 2997.300 179.760 ;
  LAYER metal3 ;
  RECT 2993.760 178.640 2997.300 179.760 ;
  LAYER metal2 ;
  RECT 2993.760 178.640 2997.300 179.760 ;
  LAYER metal1 ;
  RECT 2993.760 178.640 2997.300 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2980.120 178.640 2983.660 179.760 ;
  LAYER metal4 ;
  RECT 2980.120 178.640 2983.660 179.760 ;
  LAYER metal3 ;
  RECT 2980.120 178.640 2983.660 179.760 ;
  LAYER metal2 ;
  RECT 2980.120 178.640 2983.660 179.760 ;
  LAYER metal1 ;
  RECT 2980.120 178.640 2983.660 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2912.540 178.640 2916.080 179.760 ;
  LAYER metal4 ;
  RECT 2912.540 178.640 2916.080 179.760 ;
  LAYER metal3 ;
  RECT 2912.540 178.640 2916.080 179.760 ;
  LAYER metal2 ;
  RECT 2912.540 178.640 2916.080 179.760 ;
  LAYER metal1 ;
  RECT 2912.540 178.640 2916.080 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2899.520 178.640 2903.060 179.760 ;
  LAYER metal4 ;
  RECT 2899.520 178.640 2903.060 179.760 ;
  LAYER metal3 ;
  RECT 2899.520 178.640 2903.060 179.760 ;
  LAYER metal2 ;
  RECT 2899.520 178.640 2903.060 179.760 ;
  LAYER metal1 ;
  RECT 2899.520 178.640 2903.060 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2885.880 178.640 2889.420 179.760 ;
  LAYER metal4 ;
  RECT 2885.880 178.640 2889.420 179.760 ;
  LAYER metal3 ;
  RECT 2885.880 178.640 2889.420 179.760 ;
  LAYER metal2 ;
  RECT 2885.880 178.640 2889.420 179.760 ;
  LAYER metal1 ;
  RECT 2885.880 178.640 2889.420 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2872.240 178.640 2875.780 179.760 ;
  LAYER metal4 ;
  RECT 2872.240 178.640 2875.780 179.760 ;
  LAYER metal3 ;
  RECT 2872.240 178.640 2875.780 179.760 ;
  LAYER metal2 ;
  RECT 2872.240 178.640 2875.780 179.760 ;
  LAYER metal1 ;
  RECT 2872.240 178.640 2875.780 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2859.220 178.640 2862.760 179.760 ;
  LAYER metal4 ;
  RECT 2859.220 178.640 2862.760 179.760 ;
  LAYER metal3 ;
  RECT 2859.220 178.640 2862.760 179.760 ;
  LAYER metal2 ;
  RECT 2859.220 178.640 2862.760 179.760 ;
  LAYER metal1 ;
  RECT 2859.220 178.640 2862.760 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2845.580 178.640 2849.120 179.760 ;
  LAYER metal4 ;
  RECT 2845.580 178.640 2849.120 179.760 ;
  LAYER metal3 ;
  RECT 2845.580 178.640 2849.120 179.760 ;
  LAYER metal2 ;
  RECT 2845.580 178.640 2849.120 179.760 ;
  LAYER metal1 ;
  RECT 2845.580 178.640 2849.120 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2778.620 178.640 2782.160 179.760 ;
  LAYER metal4 ;
  RECT 2778.620 178.640 2782.160 179.760 ;
  LAYER metal3 ;
  RECT 2778.620 178.640 2782.160 179.760 ;
  LAYER metal2 ;
  RECT 2778.620 178.640 2782.160 179.760 ;
  LAYER metal1 ;
  RECT 2778.620 178.640 2782.160 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2764.980 178.640 2768.520 179.760 ;
  LAYER metal4 ;
  RECT 2764.980 178.640 2768.520 179.760 ;
  LAYER metal3 ;
  RECT 2764.980 178.640 2768.520 179.760 ;
  LAYER metal2 ;
  RECT 2764.980 178.640 2768.520 179.760 ;
  LAYER metal1 ;
  RECT 2764.980 178.640 2768.520 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2751.340 178.640 2754.880 179.760 ;
  LAYER metal4 ;
  RECT 2751.340 178.640 2754.880 179.760 ;
  LAYER metal3 ;
  RECT 2751.340 178.640 2754.880 179.760 ;
  LAYER metal2 ;
  RECT 2751.340 178.640 2754.880 179.760 ;
  LAYER metal1 ;
  RECT 2751.340 178.640 2754.880 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2738.320 178.640 2741.860 179.760 ;
  LAYER metal4 ;
  RECT 2738.320 178.640 2741.860 179.760 ;
  LAYER metal3 ;
  RECT 2738.320 178.640 2741.860 179.760 ;
  LAYER metal2 ;
  RECT 2738.320 178.640 2741.860 179.760 ;
  LAYER metal1 ;
  RECT 2738.320 178.640 2741.860 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2724.680 178.640 2728.220 179.760 ;
  LAYER metal4 ;
  RECT 2724.680 178.640 2728.220 179.760 ;
  LAYER metal3 ;
  RECT 2724.680 178.640 2728.220 179.760 ;
  LAYER metal2 ;
  RECT 2724.680 178.640 2728.220 179.760 ;
  LAYER metal1 ;
  RECT 2724.680 178.640 2728.220 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2711.040 178.640 2714.580 179.760 ;
  LAYER metal4 ;
  RECT 2711.040 178.640 2714.580 179.760 ;
  LAYER metal3 ;
  RECT 2711.040 178.640 2714.580 179.760 ;
  LAYER metal2 ;
  RECT 2711.040 178.640 2714.580 179.760 ;
  LAYER metal1 ;
  RECT 2711.040 178.640 2714.580 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2644.080 178.640 2647.620 179.760 ;
  LAYER metal4 ;
  RECT 2644.080 178.640 2647.620 179.760 ;
  LAYER metal3 ;
  RECT 2644.080 178.640 2647.620 179.760 ;
  LAYER metal2 ;
  RECT 2644.080 178.640 2647.620 179.760 ;
  LAYER metal1 ;
  RECT 2644.080 178.640 2647.620 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2630.440 178.640 2633.980 179.760 ;
  LAYER metal4 ;
  RECT 2630.440 178.640 2633.980 179.760 ;
  LAYER metal3 ;
  RECT 2630.440 178.640 2633.980 179.760 ;
  LAYER metal2 ;
  RECT 2630.440 178.640 2633.980 179.760 ;
  LAYER metal1 ;
  RECT 2630.440 178.640 2633.980 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2617.420 178.640 2620.960 179.760 ;
  LAYER metal4 ;
  RECT 2617.420 178.640 2620.960 179.760 ;
  LAYER metal3 ;
  RECT 2617.420 178.640 2620.960 179.760 ;
  LAYER metal2 ;
  RECT 2617.420 178.640 2620.960 179.760 ;
  LAYER metal1 ;
  RECT 2617.420 178.640 2620.960 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2603.780 178.640 2607.320 179.760 ;
  LAYER metal4 ;
  RECT 2603.780 178.640 2607.320 179.760 ;
  LAYER metal3 ;
  RECT 2603.780 178.640 2607.320 179.760 ;
  LAYER metal2 ;
  RECT 2603.780 178.640 2607.320 179.760 ;
  LAYER metal1 ;
  RECT 2603.780 178.640 2607.320 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2590.140 178.640 2593.680 179.760 ;
  LAYER metal4 ;
  RECT 2590.140 178.640 2593.680 179.760 ;
  LAYER metal3 ;
  RECT 2590.140 178.640 2593.680 179.760 ;
  LAYER metal2 ;
  RECT 2590.140 178.640 2593.680 179.760 ;
  LAYER metal1 ;
  RECT 2590.140 178.640 2593.680 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2577.120 178.640 2580.660 179.760 ;
  LAYER metal4 ;
  RECT 2577.120 178.640 2580.660 179.760 ;
  LAYER metal3 ;
  RECT 2577.120 178.640 2580.660 179.760 ;
  LAYER metal2 ;
  RECT 2577.120 178.640 2580.660 179.760 ;
  LAYER metal1 ;
  RECT 2577.120 178.640 2580.660 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2509.540 178.640 2513.080 179.760 ;
  LAYER metal4 ;
  RECT 2509.540 178.640 2513.080 179.760 ;
  LAYER metal3 ;
  RECT 2509.540 178.640 2513.080 179.760 ;
  LAYER metal2 ;
  RECT 2509.540 178.640 2513.080 179.760 ;
  LAYER metal1 ;
  RECT 2509.540 178.640 2513.080 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2495.900 178.640 2499.440 179.760 ;
  LAYER metal4 ;
  RECT 2495.900 178.640 2499.440 179.760 ;
  LAYER metal3 ;
  RECT 2495.900 178.640 2499.440 179.760 ;
  LAYER metal2 ;
  RECT 2495.900 178.640 2499.440 179.760 ;
  LAYER metal1 ;
  RECT 2495.900 178.640 2499.440 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2482.880 178.640 2486.420 179.760 ;
  LAYER metal4 ;
  RECT 2482.880 178.640 2486.420 179.760 ;
  LAYER metal3 ;
  RECT 2482.880 178.640 2486.420 179.760 ;
  LAYER metal2 ;
  RECT 2482.880 178.640 2486.420 179.760 ;
  LAYER metal1 ;
  RECT 2482.880 178.640 2486.420 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2469.240 178.640 2472.780 179.760 ;
  LAYER metal4 ;
  RECT 2469.240 178.640 2472.780 179.760 ;
  LAYER metal3 ;
  RECT 2469.240 178.640 2472.780 179.760 ;
  LAYER metal2 ;
  RECT 2469.240 178.640 2472.780 179.760 ;
  LAYER metal1 ;
  RECT 2469.240 178.640 2472.780 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2455.600 178.640 2459.140 179.760 ;
  LAYER metal4 ;
  RECT 2455.600 178.640 2459.140 179.760 ;
  LAYER metal3 ;
  RECT 2455.600 178.640 2459.140 179.760 ;
  LAYER metal2 ;
  RECT 2455.600 178.640 2459.140 179.760 ;
  LAYER metal1 ;
  RECT 2455.600 178.640 2459.140 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2442.580 178.640 2446.120 179.760 ;
  LAYER metal4 ;
  RECT 2442.580 178.640 2446.120 179.760 ;
  LAYER metal3 ;
  RECT 2442.580 178.640 2446.120 179.760 ;
  LAYER metal2 ;
  RECT 2442.580 178.640 2446.120 179.760 ;
  LAYER metal1 ;
  RECT 2442.580 178.640 2446.120 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2375.000 178.640 2378.540 179.760 ;
  LAYER metal4 ;
  RECT 2375.000 178.640 2378.540 179.760 ;
  LAYER metal3 ;
  RECT 2375.000 178.640 2378.540 179.760 ;
  LAYER metal2 ;
  RECT 2375.000 178.640 2378.540 179.760 ;
  LAYER metal1 ;
  RECT 2375.000 178.640 2378.540 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2361.980 178.640 2365.520 179.760 ;
  LAYER metal4 ;
  RECT 2361.980 178.640 2365.520 179.760 ;
  LAYER metal3 ;
  RECT 2361.980 178.640 2365.520 179.760 ;
  LAYER metal2 ;
  RECT 2361.980 178.640 2365.520 179.760 ;
  LAYER metal1 ;
  RECT 2361.980 178.640 2365.520 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2348.340 178.640 2351.880 179.760 ;
  LAYER metal4 ;
  RECT 2348.340 178.640 2351.880 179.760 ;
  LAYER metal3 ;
  RECT 2348.340 178.640 2351.880 179.760 ;
  LAYER metal2 ;
  RECT 2348.340 178.640 2351.880 179.760 ;
  LAYER metal1 ;
  RECT 2348.340 178.640 2351.880 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2334.700 178.640 2338.240 179.760 ;
  LAYER metal4 ;
  RECT 2334.700 178.640 2338.240 179.760 ;
  LAYER metal3 ;
  RECT 2334.700 178.640 2338.240 179.760 ;
  LAYER metal2 ;
  RECT 2334.700 178.640 2338.240 179.760 ;
  LAYER metal1 ;
  RECT 2334.700 178.640 2338.240 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2321.680 178.640 2325.220 179.760 ;
  LAYER metal4 ;
  RECT 2321.680 178.640 2325.220 179.760 ;
  LAYER metal3 ;
  RECT 2321.680 178.640 2325.220 179.760 ;
  LAYER metal2 ;
  RECT 2321.680 178.640 2325.220 179.760 ;
  LAYER metal1 ;
  RECT 2321.680 178.640 2325.220 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2308.040 178.640 2311.580 179.760 ;
  LAYER metal4 ;
  RECT 2308.040 178.640 2311.580 179.760 ;
  LAYER metal3 ;
  RECT 2308.040 178.640 2311.580 179.760 ;
  LAYER metal2 ;
  RECT 2308.040 178.640 2311.580 179.760 ;
  LAYER metal1 ;
  RECT 2308.040 178.640 2311.580 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2241.080 178.640 2244.620 179.760 ;
  LAYER metal4 ;
  RECT 2241.080 178.640 2244.620 179.760 ;
  LAYER metal3 ;
  RECT 2241.080 178.640 2244.620 179.760 ;
  LAYER metal2 ;
  RECT 2241.080 178.640 2244.620 179.760 ;
  LAYER metal1 ;
  RECT 2241.080 178.640 2244.620 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2227.440 178.640 2230.980 179.760 ;
  LAYER metal4 ;
  RECT 2227.440 178.640 2230.980 179.760 ;
  LAYER metal3 ;
  RECT 2227.440 178.640 2230.980 179.760 ;
  LAYER metal2 ;
  RECT 2227.440 178.640 2230.980 179.760 ;
  LAYER metal1 ;
  RECT 2227.440 178.640 2230.980 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2213.800 178.640 2217.340 179.760 ;
  LAYER metal4 ;
  RECT 2213.800 178.640 2217.340 179.760 ;
  LAYER metal3 ;
  RECT 2213.800 178.640 2217.340 179.760 ;
  LAYER metal2 ;
  RECT 2213.800 178.640 2217.340 179.760 ;
  LAYER metal1 ;
  RECT 2213.800 178.640 2217.340 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2200.780 178.640 2204.320 179.760 ;
  LAYER metal4 ;
  RECT 2200.780 178.640 2204.320 179.760 ;
  LAYER metal3 ;
  RECT 2200.780 178.640 2204.320 179.760 ;
  LAYER metal2 ;
  RECT 2200.780 178.640 2204.320 179.760 ;
  LAYER metal1 ;
  RECT 2200.780 178.640 2204.320 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2187.140 178.640 2190.680 179.760 ;
  LAYER metal4 ;
  RECT 2187.140 178.640 2190.680 179.760 ;
  LAYER metal3 ;
  RECT 2187.140 178.640 2190.680 179.760 ;
  LAYER metal2 ;
  RECT 2187.140 178.640 2190.680 179.760 ;
  LAYER metal1 ;
  RECT 2187.140 178.640 2190.680 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2173.500 178.640 2177.040 179.760 ;
  LAYER metal4 ;
  RECT 2173.500 178.640 2177.040 179.760 ;
  LAYER metal3 ;
  RECT 2173.500 178.640 2177.040 179.760 ;
  LAYER metal2 ;
  RECT 2173.500 178.640 2177.040 179.760 ;
  LAYER metal1 ;
  RECT 2173.500 178.640 2177.040 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2106.540 178.640 2110.080 179.760 ;
  LAYER metal4 ;
  RECT 2106.540 178.640 2110.080 179.760 ;
  LAYER metal3 ;
  RECT 2106.540 178.640 2110.080 179.760 ;
  LAYER metal2 ;
  RECT 2106.540 178.640 2110.080 179.760 ;
  LAYER metal1 ;
  RECT 2106.540 178.640 2110.080 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2092.900 178.640 2096.440 179.760 ;
  LAYER metal4 ;
  RECT 2092.900 178.640 2096.440 179.760 ;
  LAYER metal3 ;
  RECT 2092.900 178.640 2096.440 179.760 ;
  LAYER metal2 ;
  RECT 2092.900 178.640 2096.440 179.760 ;
  LAYER metal1 ;
  RECT 2092.900 178.640 2096.440 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2079.260 178.640 2082.800 179.760 ;
  LAYER metal4 ;
  RECT 2079.260 178.640 2082.800 179.760 ;
  LAYER metal3 ;
  RECT 2079.260 178.640 2082.800 179.760 ;
  LAYER metal2 ;
  RECT 2079.260 178.640 2082.800 179.760 ;
  LAYER metal1 ;
  RECT 2079.260 178.640 2082.800 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2066.240 178.640 2069.780 179.760 ;
  LAYER metal4 ;
  RECT 2066.240 178.640 2069.780 179.760 ;
  LAYER metal3 ;
  RECT 2066.240 178.640 2069.780 179.760 ;
  LAYER metal2 ;
  RECT 2066.240 178.640 2069.780 179.760 ;
  LAYER metal1 ;
  RECT 2066.240 178.640 2069.780 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2052.600 178.640 2056.140 179.760 ;
  LAYER metal4 ;
  RECT 2052.600 178.640 2056.140 179.760 ;
  LAYER metal3 ;
  RECT 2052.600 178.640 2056.140 179.760 ;
  LAYER metal2 ;
  RECT 2052.600 178.640 2056.140 179.760 ;
  LAYER metal1 ;
  RECT 2052.600 178.640 2056.140 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2038.960 178.640 2042.500 179.760 ;
  LAYER metal4 ;
  RECT 2038.960 178.640 2042.500 179.760 ;
  LAYER metal3 ;
  RECT 2038.960 178.640 2042.500 179.760 ;
  LAYER metal2 ;
  RECT 2038.960 178.640 2042.500 179.760 ;
  LAYER metal1 ;
  RECT 2038.960 178.640 2042.500 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1972.000 178.640 1975.540 179.760 ;
  LAYER metal4 ;
  RECT 1972.000 178.640 1975.540 179.760 ;
  LAYER metal3 ;
  RECT 1972.000 178.640 1975.540 179.760 ;
  LAYER metal2 ;
  RECT 1972.000 178.640 1975.540 179.760 ;
  LAYER metal1 ;
  RECT 1972.000 178.640 1975.540 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1958.360 178.640 1961.900 179.760 ;
  LAYER metal4 ;
  RECT 1958.360 178.640 1961.900 179.760 ;
  LAYER metal3 ;
  RECT 1958.360 178.640 1961.900 179.760 ;
  LAYER metal2 ;
  RECT 1958.360 178.640 1961.900 179.760 ;
  LAYER metal1 ;
  RECT 1958.360 178.640 1961.900 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1945.340 178.640 1948.880 179.760 ;
  LAYER metal4 ;
  RECT 1945.340 178.640 1948.880 179.760 ;
  LAYER metal3 ;
  RECT 1945.340 178.640 1948.880 179.760 ;
  LAYER metal2 ;
  RECT 1945.340 178.640 1948.880 179.760 ;
  LAYER metal1 ;
  RECT 1945.340 178.640 1948.880 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1931.700 178.640 1935.240 179.760 ;
  LAYER metal4 ;
  RECT 1931.700 178.640 1935.240 179.760 ;
  LAYER metal3 ;
  RECT 1931.700 178.640 1935.240 179.760 ;
  LAYER metal2 ;
  RECT 1931.700 178.640 1935.240 179.760 ;
  LAYER metal1 ;
  RECT 1931.700 178.640 1935.240 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1918.060 178.640 1921.600 179.760 ;
  LAYER metal4 ;
  RECT 1918.060 178.640 1921.600 179.760 ;
  LAYER metal3 ;
  RECT 1918.060 178.640 1921.600 179.760 ;
  LAYER metal2 ;
  RECT 1918.060 178.640 1921.600 179.760 ;
  LAYER metal1 ;
  RECT 1918.060 178.640 1921.600 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1905.040 178.640 1908.580 179.760 ;
  LAYER metal4 ;
  RECT 1905.040 178.640 1908.580 179.760 ;
  LAYER metal3 ;
  RECT 1905.040 178.640 1908.580 179.760 ;
  LAYER metal2 ;
  RECT 1905.040 178.640 1908.580 179.760 ;
  LAYER metal1 ;
  RECT 1905.040 178.640 1908.580 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1837.460 178.640 1841.000 179.760 ;
  LAYER metal4 ;
  RECT 1837.460 178.640 1841.000 179.760 ;
  LAYER metal3 ;
  RECT 1837.460 178.640 1841.000 179.760 ;
  LAYER metal2 ;
  RECT 1837.460 178.640 1841.000 179.760 ;
  LAYER metal1 ;
  RECT 1837.460 178.640 1841.000 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1826.300 178.640 1829.840 179.760 ;
  LAYER metal4 ;
  RECT 1826.300 178.640 1829.840 179.760 ;
  LAYER metal3 ;
  RECT 1826.300 178.640 1829.840 179.760 ;
  LAYER metal2 ;
  RECT 1826.300 178.640 1829.840 179.760 ;
  LAYER metal1 ;
  RECT 1826.300 178.640 1829.840 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1810.180 178.640 1813.720 179.760 ;
  LAYER metal4 ;
  RECT 1810.180 178.640 1813.720 179.760 ;
  LAYER metal3 ;
  RECT 1810.180 178.640 1813.720 179.760 ;
  LAYER metal2 ;
  RECT 1810.180 178.640 1813.720 179.760 ;
  LAYER metal1 ;
  RECT 1810.180 178.640 1813.720 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1801.500 178.640 1805.040 179.760 ;
  LAYER metal4 ;
  RECT 1801.500 178.640 1805.040 179.760 ;
  LAYER metal3 ;
  RECT 1801.500 178.640 1805.040 179.760 ;
  LAYER metal2 ;
  RECT 1801.500 178.640 1805.040 179.760 ;
  LAYER metal1 ;
  RECT 1801.500 178.640 1805.040 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1792.820 178.640 1796.360 179.760 ;
  LAYER metal4 ;
  RECT 1792.820 178.640 1796.360 179.760 ;
  LAYER metal3 ;
  RECT 1792.820 178.640 1796.360 179.760 ;
  LAYER metal2 ;
  RECT 1792.820 178.640 1796.360 179.760 ;
  LAYER metal1 ;
  RECT 1792.820 178.640 1796.360 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1779.800 178.640 1783.340 179.760 ;
  LAYER metal4 ;
  RECT 1779.800 178.640 1783.340 179.760 ;
  LAYER metal3 ;
  RECT 1779.800 178.640 1783.340 179.760 ;
  LAYER metal2 ;
  RECT 1779.800 178.640 1783.340 179.760 ;
  LAYER metal1 ;
  RECT 1779.800 178.640 1783.340 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1694.860 178.640 1698.400 179.760 ;
  LAYER metal4 ;
  RECT 1694.860 178.640 1698.400 179.760 ;
  LAYER metal3 ;
  RECT 1694.860 178.640 1698.400 179.760 ;
  LAYER metal2 ;
  RECT 1694.860 178.640 1698.400 179.760 ;
  LAYER metal1 ;
  RECT 1694.860 178.640 1698.400 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1681.220 178.640 1684.760 179.760 ;
  LAYER metal4 ;
  RECT 1681.220 178.640 1684.760 179.760 ;
  LAYER metal3 ;
  RECT 1681.220 178.640 1684.760 179.760 ;
  LAYER metal2 ;
  RECT 1681.220 178.640 1684.760 179.760 ;
  LAYER metal1 ;
  RECT 1681.220 178.640 1684.760 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1668.200 178.640 1671.740 179.760 ;
  LAYER metal4 ;
  RECT 1668.200 178.640 1671.740 179.760 ;
  LAYER metal3 ;
  RECT 1668.200 178.640 1671.740 179.760 ;
  LAYER metal2 ;
  RECT 1668.200 178.640 1671.740 179.760 ;
  LAYER metal1 ;
  RECT 1668.200 178.640 1671.740 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1654.560 178.640 1658.100 179.760 ;
  LAYER metal4 ;
  RECT 1654.560 178.640 1658.100 179.760 ;
  LAYER metal3 ;
  RECT 1654.560 178.640 1658.100 179.760 ;
  LAYER metal2 ;
  RECT 1654.560 178.640 1658.100 179.760 ;
  LAYER metal1 ;
  RECT 1654.560 178.640 1658.100 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1640.920 178.640 1644.460 179.760 ;
  LAYER metal4 ;
  RECT 1640.920 178.640 1644.460 179.760 ;
  LAYER metal3 ;
  RECT 1640.920 178.640 1644.460 179.760 ;
  LAYER metal2 ;
  RECT 1640.920 178.640 1644.460 179.760 ;
  LAYER metal1 ;
  RECT 1640.920 178.640 1644.460 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1627.900 178.640 1631.440 179.760 ;
  LAYER metal4 ;
  RECT 1627.900 178.640 1631.440 179.760 ;
  LAYER metal3 ;
  RECT 1627.900 178.640 1631.440 179.760 ;
  LAYER metal2 ;
  RECT 1627.900 178.640 1631.440 179.760 ;
  LAYER metal1 ;
  RECT 1627.900 178.640 1631.440 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1560.320 178.640 1563.860 179.760 ;
  LAYER metal4 ;
  RECT 1560.320 178.640 1563.860 179.760 ;
  LAYER metal3 ;
  RECT 1560.320 178.640 1563.860 179.760 ;
  LAYER metal2 ;
  RECT 1560.320 178.640 1563.860 179.760 ;
  LAYER metal1 ;
  RECT 1560.320 178.640 1563.860 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1547.300 178.640 1550.840 179.760 ;
  LAYER metal4 ;
  RECT 1547.300 178.640 1550.840 179.760 ;
  LAYER metal3 ;
  RECT 1547.300 178.640 1550.840 179.760 ;
  LAYER metal2 ;
  RECT 1547.300 178.640 1550.840 179.760 ;
  LAYER metal1 ;
  RECT 1547.300 178.640 1550.840 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1533.660 178.640 1537.200 179.760 ;
  LAYER metal4 ;
  RECT 1533.660 178.640 1537.200 179.760 ;
  LAYER metal3 ;
  RECT 1533.660 178.640 1537.200 179.760 ;
  LAYER metal2 ;
  RECT 1533.660 178.640 1537.200 179.760 ;
  LAYER metal1 ;
  RECT 1533.660 178.640 1537.200 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1520.020 178.640 1523.560 179.760 ;
  LAYER metal4 ;
  RECT 1520.020 178.640 1523.560 179.760 ;
  LAYER metal3 ;
  RECT 1520.020 178.640 1523.560 179.760 ;
  LAYER metal2 ;
  RECT 1520.020 178.640 1523.560 179.760 ;
  LAYER metal1 ;
  RECT 1520.020 178.640 1523.560 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1507.000 178.640 1510.540 179.760 ;
  LAYER metal4 ;
  RECT 1507.000 178.640 1510.540 179.760 ;
  LAYER metal3 ;
  RECT 1507.000 178.640 1510.540 179.760 ;
  LAYER metal2 ;
  RECT 1507.000 178.640 1510.540 179.760 ;
  LAYER metal1 ;
  RECT 1507.000 178.640 1510.540 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1493.360 178.640 1496.900 179.760 ;
  LAYER metal4 ;
  RECT 1493.360 178.640 1496.900 179.760 ;
  LAYER metal3 ;
  RECT 1493.360 178.640 1496.900 179.760 ;
  LAYER metal2 ;
  RECT 1493.360 178.640 1496.900 179.760 ;
  LAYER metal1 ;
  RECT 1493.360 178.640 1496.900 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1426.400 178.640 1429.940 179.760 ;
  LAYER metal4 ;
  RECT 1426.400 178.640 1429.940 179.760 ;
  LAYER metal3 ;
  RECT 1426.400 178.640 1429.940 179.760 ;
  LAYER metal2 ;
  RECT 1426.400 178.640 1429.940 179.760 ;
  LAYER metal1 ;
  RECT 1426.400 178.640 1429.940 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1412.760 178.640 1416.300 179.760 ;
  LAYER metal4 ;
  RECT 1412.760 178.640 1416.300 179.760 ;
  LAYER metal3 ;
  RECT 1412.760 178.640 1416.300 179.760 ;
  LAYER metal2 ;
  RECT 1412.760 178.640 1416.300 179.760 ;
  LAYER metal1 ;
  RECT 1412.760 178.640 1416.300 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1399.120 178.640 1402.660 179.760 ;
  LAYER metal4 ;
  RECT 1399.120 178.640 1402.660 179.760 ;
  LAYER metal3 ;
  RECT 1399.120 178.640 1402.660 179.760 ;
  LAYER metal2 ;
  RECT 1399.120 178.640 1402.660 179.760 ;
  LAYER metal1 ;
  RECT 1399.120 178.640 1402.660 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1386.100 178.640 1389.640 179.760 ;
  LAYER metal4 ;
  RECT 1386.100 178.640 1389.640 179.760 ;
  LAYER metal3 ;
  RECT 1386.100 178.640 1389.640 179.760 ;
  LAYER metal2 ;
  RECT 1386.100 178.640 1389.640 179.760 ;
  LAYER metal1 ;
  RECT 1386.100 178.640 1389.640 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1372.460 178.640 1376.000 179.760 ;
  LAYER metal4 ;
  RECT 1372.460 178.640 1376.000 179.760 ;
  LAYER metal3 ;
  RECT 1372.460 178.640 1376.000 179.760 ;
  LAYER metal2 ;
  RECT 1372.460 178.640 1376.000 179.760 ;
  LAYER metal1 ;
  RECT 1372.460 178.640 1376.000 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1358.820 178.640 1362.360 179.760 ;
  LAYER metal4 ;
  RECT 1358.820 178.640 1362.360 179.760 ;
  LAYER metal3 ;
  RECT 1358.820 178.640 1362.360 179.760 ;
  LAYER metal2 ;
  RECT 1358.820 178.640 1362.360 179.760 ;
  LAYER metal1 ;
  RECT 1358.820 178.640 1362.360 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1291.860 178.640 1295.400 179.760 ;
  LAYER metal4 ;
  RECT 1291.860 178.640 1295.400 179.760 ;
  LAYER metal3 ;
  RECT 1291.860 178.640 1295.400 179.760 ;
  LAYER metal2 ;
  RECT 1291.860 178.640 1295.400 179.760 ;
  LAYER metal1 ;
  RECT 1291.860 178.640 1295.400 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1278.220 178.640 1281.760 179.760 ;
  LAYER metal4 ;
  RECT 1278.220 178.640 1281.760 179.760 ;
  LAYER metal3 ;
  RECT 1278.220 178.640 1281.760 179.760 ;
  LAYER metal2 ;
  RECT 1278.220 178.640 1281.760 179.760 ;
  LAYER metal1 ;
  RECT 1278.220 178.640 1281.760 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1264.580 178.640 1268.120 179.760 ;
  LAYER metal4 ;
  RECT 1264.580 178.640 1268.120 179.760 ;
  LAYER metal3 ;
  RECT 1264.580 178.640 1268.120 179.760 ;
  LAYER metal2 ;
  RECT 1264.580 178.640 1268.120 179.760 ;
  LAYER metal1 ;
  RECT 1264.580 178.640 1268.120 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1251.560 178.640 1255.100 179.760 ;
  LAYER metal4 ;
  RECT 1251.560 178.640 1255.100 179.760 ;
  LAYER metal3 ;
  RECT 1251.560 178.640 1255.100 179.760 ;
  LAYER metal2 ;
  RECT 1251.560 178.640 1255.100 179.760 ;
  LAYER metal1 ;
  RECT 1251.560 178.640 1255.100 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1237.920 178.640 1241.460 179.760 ;
  LAYER metal4 ;
  RECT 1237.920 178.640 1241.460 179.760 ;
  LAYER metal3 ;
  RECT 1237.920 178.640 1241.460 179.760 ;
  LAYER metal2 ;
  RECT 1237.920 178.640 1241.460 179.760 ;
  LAYER metal1 ;
  RECT 1237.920 178.640 1241.460 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1224.280 178.640 1227.820 179.760 ;
  LAYER metal4 ;
  RECT 1224.280 178.640 1227.820 179.760 ;
  LAYER metal3 ;
  RECT 1224.280 178.640 1227.820 179.760 ;
  LAYER metal2 ;
  RECT 1224.280 178.640 1227.820 179.760 ;
  LAYER metal1 ;
  RECT 1224.280 178.640 1227.820 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1157.320 178.640 1160.860 179.760 ;
  LAYER metal4 ;
  RECT 1157.320 178.640 1160.860 179.760 ;
  LAYER metal3 ;
  RECT 1157.320 178.640 1160.860 179.760 ;
  LAYER metal2 ;
  RECT 1157.320 178.640 1160.860 179.760 ;
  LAYER metal1 ;
  RECT 1157.320 178.640 1160.860 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1143.680 178.640 1147.220 179.760 ;
  LAYER metal4 ;
  RECT 1143.680 178.640 1147.220 179.760 ;
  LAYER metal3 ;
  RECT 1143.680 178.640 1147.220 179.760 ;
  LAYER metal2 ;
  RECT 1143.680 178.640 1147.220 179.760 ;
  LAYER metal1 ;
  RECT 1143.680 178.640 1147.220 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1130.660 178.640 1134.200 179.760 ;
  LAYER metal4 ;
  RECT 1130.660 178.640 1134.200 179.760 ;
  LAYER metal3 ;
  RECT 1130.660 178.640 1134.200 179.760 ;
  LAYER metal2 ;
  RECT 1130.660 178.640 1134.200 179.760 ;
  LAYER metal1 ;
  RECT 1130.660 178.640 1134.200 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1117.020 178.640 1120.560 179.760 ;
  LAYER metal4 ;
  RECT 1117.020 178.640 1120.560 179.760 ;
  LAYER metal3 ;
  RECT 1117.020 178.640 1120.560 179.760 ;
  LAYER metal2 ;
  RECT 1117.020 178.640 1120.560 179.760 ;
  LAYER metal1 ;
  RECT 1117.020 178.640 1120.560 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1103.380 178.640 1106.920 179.760 ;
  LAYER metal4 ;
  RECT 1103.380 178.640 1106.920 179.760 ;
  LAYER metal3 ;
  RECT 1103.380 178.640 1106.920 179.760 ;
  LAYER metal2 ;
  RECT 1103.380 178.640 1106.920 179.760 ;
  LAYER metal1 ;
  RECT 1103.380 178.640 1106.920 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1090.360 178.640 1093.900 179.760 ;
  LAYER metal4 ;
  RECT 1090.360 178.640 1093.900 179.760 ;
  LAYER metal3 ;
  RECT 1090.360 178.640 1093.900 179.760 ;
  LAYER metal2 ;
  RECT 1090.360 178.640 1093.900 179.760 ;
  LAYER metal1 ;
  RECT 1090.360 178.640 1093.900 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1022.780 178.640 1026.320 179.760 ;
  LAYER metal4 ;
  RECT 1022.780 178.640 1026.320 179.760 ;
  LAYER metal3 ;
  RECT 1022.780 178.640 1026.320 179.760 ;
  LAYER metal2 ;
  RECT 1022.780 178.640 1026.320 179.760 ;
  LAYER metal1 ;
  RECT 1022.780 178.640 1026.320 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1009.760 178.640 1013.300 179.760 ;
  LAYER metal4 ;
  RECT 1009.760 178.640 1013.300 179.760 ;
  LAYER metal3 ;
  RECT 1009.760 178.640 1013.300 179.760 ;
  LAYER metal2 ;
  RECT 1009.760 178.640 1013.300 179.760 ;
  LAYER metal1 ;
  RECT 1009.760 178.640 1013.300 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 996.120 178.640 999.660 179.760 ;
  LAYER metal4 ;
  RECT 996.120 178.640 999.660 179.760 ;
  LAYER metal3 ;
  RECT 996.120 178.640 999.660 179.760 ;
  LAYER metal2 ;
  RECT 996.120 178.640 999.660 179.760 ;
  LAYER metal1 ;
  RECT 996.120 178.640 999.660 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 982.480 178.640 986.020 179.760 ;
  LAYER metal4 ;
  RECT 982.480 178.640 986.020 179.760 ;
  LAYER metal3 ;
  RECT 982.480 178.640 986.020 179.760 ;
  LAYER metal2 ;
  RECT 982.480 178.640 986.020 179.760 ;
  LAYER metal1 ;
  RECT 982.480 178.640 986.020 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 969.460 178.640 973.000 179.760 ;
  LAYER metal4 ;
  RECT 969.460 178.640 973.000 179.760 ;
  LAYER metal3 ;
  RECT 969.460 178.640 973.000 179.760 ;
  LAYER metal2 ;
  RECT 969.460 178.640 973.000 179.760 ;
  LAYER metal1 ;
  RECT 969.460 178.640 973.000 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 955.820 178.640 959.360 179.760 ;
  LAYER metal4 ;
  RECT 955.820 178.640 959.360 179.760 ;
  LAYER metal3 ;
  RECT 955.820 178.640 959.360 179.760 ;
  LAYER metal2 ;
  RECT 955.820 178.640 959.360 179.760 ;
  LAYER metal1 ;
  RECT 955.820 178.640 959.360 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 888.240 178.640 891.780 179.760 ;
  LAYER metal4 ;
  RECT 888.240 178.640 891.780 179.760 ;
  LAYER metal3 ;
  RECT 888.240 178.640 891.780 179.760 ;
  LAYER metal2 ;
  RECT 888.240 178.640 891.780 179.760 ;
  LAYER metal1 ;
  RECT 888.240 178.640 891.780 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 877.080 178.640 880.620 179.760 ;
  LAYER metal4 ;
  RECT 877.080 178.640 880.620 179.760 ;
  LAYER metal3 ;
  RECT 877.080 178.640 880.620 179.760 ;
  LAYER metal2 ;
  RECT 877.080 178.640 880.620 179.760 ;
  LAYER metal1 ;
  RECT 877.080 178.640 880.620 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 861.580 178.640 865.120 179.760 ;
  LAYER metal4 ;
  RECT 861.580 178.640 865.120 179.760 ;
  LAYER metal3 ;
  RECT 861.580 178.640 865.120 179.760 ;
  LAYER metal2 ;
  RECT 861.580 178.640 865.120 179.760 ;
  LAYER metal1 ;
  RECT 861.580 178.640 865.120 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 847.940 178.640 851.480 179.760 ;
  LAYER metal4 ;
  RECT 847.940 178.640 851.480 179.760 ;
  LAYER metal3 ;
  RECT 847.940 178.640 851.480 179.760 ;
  LAYER metal2 ;
  RECT 847.940 178.640 851.480 179.760 ;
  LAYER metal1 ;
  RECT 847.940 178.640 851.480 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 834.920 178.640 838.460 179.760 ;
  LAYER metal4 ;
  RECT 834.920 178.640 838.460 179.760 ;
  LAYER metal3 ;
  RECT 834.920 178.640 838.460 179.760 ;
  LAYER metal2 ;
  RECT 834.920 178.640 838.460 179.760 ;
  LAYER metal1 ;
  RECT 834.920 178.640 838.460 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 821.280 178.640 824.820 179.760 ;
  LAYER metal4 ;
  RECT 821.280 178.640 824.820 179.760 ;
  LAYER metal3 ;
  RECT 821.280 178.640 824.820 179.760 ;
  LAYER metal2 ;
  RECT 821.280 178.640 824.820 179.760 ;
  LAYER metal1 ;
  RECT 821.280 178.640 824.820 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 754.320 178.640 757.860 179.760 ;
  LAYER metal4 ;
  RECT 754.320 178.640 757.860 179.760 ;
  LAYER metal3 ;
  RECT 754.320 178.640 757.860 179.760 ;
  LAYER metal2 ;
  RECT 754.320 178.640 757.860 179.760 ;
  LAYER metal1 ;
  RECT 754.320 178.640 757.860 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 740.680 178.640 744.220 179.760 ;
  LAYER metal4 ;
  RECT 740.680 178.640 744.220 179.760 ;
  LAYER metal3 ;
  RECT 740.680 178.640 744.220 179.760 ;
  LAYER metal2 ;
  RECT 740.680 178.640 744.220 179.760 ;
  LAYER metal1 ;
  RECT 740.680 178.640 744.220 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 727.040 178.640 730.580 179.760 ;
  LAYER metal4 ;
  RECT 727.040 178.640 730.580 179.760 ;
  LAYER metal3 ;
  RECT 727.040 178.640 730.580 179.760 ;
  LAYER metal2 ;
  RECT 727.040 178.640 730.580 179.760 ;
  LAYER metal1 ;
  RECT 727.040 178.640 730.580 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 714.020 178.640 717.560 179.760 ;
  LAYER metal4 ;
  RECT 714.020 178.640 717.560 179.760 ;
  LAYER metal3 ;
  RECT 714.020 178.640 717.560 179.760 ;
  LAYER metal2 ;
  RECT 714.020 178.640 717.560 179.760 ;
  LAYER metal1 ;
  RECT 714.020 178.640 717.560 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 700.380 178.640 703.920 179.760 ;
  LAYER metal4 ;
  RECT 700.380 178.640 703.920 179.760 ;
  LAYER metal3 ;
  RECT 700.380 178.640 703.920 179.760 ;
  LAYER metal2 ;
  RECT 700.380 178.640 703.920 179.760 ;
  LAYER metal1 ;
  RECT 700.380 178.640 703.920 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 686.740 178.640 690.280 179.760 ;
  LAYER metal4 ;
  RECT 686.740 178.640 690.280 179.760 ;
  LAYER metal3 ;
  RECT 686.740 178.640 690.280 179.760 ;
  LAYER metal2 ;
  RECT 686.740 178.640 690.280 179.760 ;
  LAYER metal1 ;
  RECT 686.740 178.640 690.280 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 619.780 178.640 623.320 179.760 ;
  LAYER metal4 ;
  RECT 619.780 178.640 623.320 179.760 ;
  LAYER metal3 ;
  RECT 619.780 178.640 623.320 179.760 ;
  LAYER metal2 ;
  RECT 619.780 178.640 623.320 179.760 ;
  LAYER metal1 ;
  RECT 619.780 178.640 623.320 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 606.140 178.640 609.680 179.760 ;
  LAYER metal4 ;
  RECT 606.140 178.640 609.680 179.760 ;
  LAYER metal3 ;
  RECT 606.140 178.640 609.680 179.760 ;
  LAYER metal2 ;
  RECT 606.140 178.640 609.680 179.760 ;
  LAYER metal1 ;
  RECT 606.140 178.640 609.680 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 593.120 178.640 596.660 179.760 ;
  LAYER metal4 ;
  RECT 593.120 178.640 596.660 179.760 ;
  LAYER metal3 ;
  RECT 593.120 178.640 596.660 179.760 ;
  LAYER metal2 ;
  RECT 593.120 178.640 596.660 179.760 ;
  LAYER metal1 ;
  RECT 593.120 178.640 596.660 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 579.480 178.640 583.020 179.760 ;
  LAYER metal4 ;
  RECT 579.480 178.640 583.020 179.760 ;
  LAYER metal3 ;
  RECT 579.480 178.640 583.020 179.760 ;
  LAYER metal2 ;
  RECT 579.480 178.640 583.020 179.760 ;
  LAYER metal1 ;
  RECT 579.480 178.640 583.020 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 565.840 178.640 569.380 179.760 ;
  LAYER metal4 ;
  RECT 565.840 178.640 569.380 179.760 ;
  LAYER metal3 ;
  RECT 565.840 178.640 569.380 179.760 ;
  LAYER metal2 ;
  RECT 565.840 178.640 569.380 179.760 ;
  LAYER metal1 ;
  RECT 565.840 178.640 569.380 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 552.820 178.640 556.360 179.760 ;
  LAYER metal4 ;
  RECT 552.820 178.640 556.360 179.760 ;
  LAYER metal3 ;
  RECT 552.820 178.640 556.360 179.760 ;
  LAYER metal2 ;
  RECT 552.820 178.640 556.360 179.760 ;
  LAYER metal1 ;
  RECT 552.820 178.640 556.360 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 485.240 178.640 488.780 179.760 ;
  LAYER metal4 ;
  RECT 485.240 178.640 488.780 179.760 ;
  LAYER metal3 ;
  RECT 485.240 178.640 488.780 179.760 ;
  LAYER metal2 ;
  RECT 485.240 178.640 488.780 179.760 ;
  LAYER metal1 ;
  RECT 485.240 178.640 488.780 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 471.600 178.640 475.140 179.760 ;
  LAYER metal4 ;
  RECT 471.600 178.640 475.140 179.760 ;
  LAYER metal3 ;
  RECT 471.600 178.640 475.140 179.760 ;
  LAYER metal2 ;
  RECT 471.600 178.640 475.140 179.760 ;
  LAYER metal1 ;
  RECT 471.600 178.640 475.140 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 458.580 178.640 462.120 179.760 ;
  LAYER metal4 ;
  RECT 458.580 178.640 462.120 179.760 ;
  LAYER metal3 ;
  RECT 458.580 178.640 462.120 179.760 ;
  LAYER metal2 ;
  RECT 458.580 178.640 462.120 179.760 ;
  LAYER metal1 ;
  RECT 458.580 178.640 462.120 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 447.420 178.640 450.960 179.760 ;
  LAYER metal4 ;
  RECT 447.420 178.640 450.960 179.760 ;
  LAYER metal3 ;
  RECT 447.420 178.640 450.960 179.760 ;
  LAYER metal2 ;
  RECT 447.420 178.640 450.960 179.760 ;
  LAYER metal1 ;
  RECT 447.420 178.640 450.960 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 431.300 178.640 434.840 179.760 ;
  LAYER metal4 ;
  RECT 431.300 178.640 434.840 179.760 ;
  LAYER metal3 ;
  RECT 431.300 178.640 434.840 179.760 ;
  LAYER metal2 ;
  RECT 431.300 178.640 434.840 179.760 ;
  LAYER metal1 ;
  RECT 431.300 178.640 434.840 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 418.280 178.640 421.820 179.760 ;
  LAYER metal4 ;
  RECT 418.280 178.640 421.820 179.760 ;
  LAYER metal3 ;
  RECT 418.280 178.640 421.820 179.760 ;
  LAYER metal2 ;
  RECT 418.280 178.640 421.820 179.760 ;
  LAYER metal1 ;
  RECT 418.280 178.640 421.820 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 350.700 178.640 354.240 179.760 ;
  LAYER metal4 ;
  RECT 350.700 178.640 354.240 179.760 ;
  LAYER metal3 ;
  RECT 350.700 178.640 354.240 179.760 ;
  LAYER metal2 ;
  RECT 350.700 178.640 354.240 179.760 ;
  LAYER metal1 ;
  RECT 350.700 178.640 354.240 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 337.680 178.640 341.220 179.760 ;
  LAYER metal4 ;
  RECT 337.680 178.640 341.220 179.760 ;
  LAYER metal3 ;
  RECT 337.680 178.640 341.220 179.760 ;
  LAYER metal2 ;
  RECT 337.680 178.640 341.220 179.760 ;
  LAYER metal1 ;
  RECT 337.680 178.640 341.220 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 324.040 178.640 327.580 179.760 ;
  LAYER metal4 ;
  RECT 324.040 178.640 327.580 179.760 ;
  LAYER metal3 ;
  RECT 324.040 178.640 327.580 179.760 ;
  LAYER metal2 ;
  RECT 324.040 178.640 327.580 179.760 ;
  LAYER metal1 ;
  RECT 324.040 178.640 327.580 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 310.400 178.640 313.940 179.760 ;
  LAYER metal4 ;
  RECT 310.400 178.640 313.940 179.760 ;
  LAYER metal3 ;
  RECT 310.400 178.640 313.940 179.760 ;
  LAYER metal2 ;
  RECT 310.400 178.640 313.940 179.760 ;
  LAYER metal1 ;
  RECT 310.400 178.640 313.940 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 297.380 178.640 300.920 179.760 ;
  LAYER metal4 ;
  RECT 297.380 178.640 300.920 179.760 ;
  LAYER metal3 ;
  RECT 297.380 178.640 300.920 179.760 ;
  LAYER metal2 ;
  RECT 297.380 178.640 300.920 179.760 ;
  LAYER metal1 ;
  RECT 297.380 178.640 300.920 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 283.740 178.640 287.280 179.760 ;
  LAYER metal4 ;
  RECT 283.740 178.640 287.280 179.760 ;
  LAYER metal3 ;
  RECT 283.740 178.640 287.280 179.760 ;
  LAYER metal2 ;
  RECT 283.740 178.640 287.280 179.760 ;
  LAYER metal1 ;
  RECT 283.740 178.640 287.280 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 216.780 178.640 220.320 179.760 ;
  LAYER metal4 ;
  RECT 216.780 178.640 220.320 179.760 ;
  LAYER metal3 ;
  RECT 216.780 178.640 220.320 179.760 ;
  LAYER metal2 ;
  RECT 216.780 178.640 220.320 179.760 ;
  LAYER metal1 ;
  RECT 216.780 178.640 220.320 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 203.140 178.640 206.680 179.760 ;
  LAYER metal4 ;
  RECT 203.140 178.640 206.680 179.760 ;
  LAYER metal3 ;
  RECT 203.140 178.640 206.680 179.760 ;
  LAYER metal2 ;
  RECT 203.140 178.640 206.680 179.760 ;
  LAYER metal1 ;
  RECT 203.140 178.640 206.680 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 189.500 178.640 193.040 179.760 ;
  LAYER metal4 ;
  RECT 189.500 178.640 193.040 179.760 ;
  LAYER metal3 ;
  RECT 189.500 178.640 193.040 179.760 ;
  LAYER metal2 ;
  RECT 189.500 178.640 193.040 179.760 ;
  LAYER metal1 ;
  RECT 189.500 178.640 193.040 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 176.480 178.640 180.020 179.760 ;
  LAYER metal4 ;
  RECT 176.480 178.640 180.020 179.760 ;
  LAYER metal3 ;
  RECT 176.480 178.640 180.020 179.760 ;
  LAYER metal2 ;
  RECT 176.480 178.640 180.020 179.760 ;
  LAYER metal1 ;
  RECT 176.480 178.640 180.020 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 162.840 178.640 166.380 179.760 ;
  LAYER metal4 ;
  RECT 162.840 178.640 166.380 179.760 ;
  LAYER metal3 ;
  RECT 162.840 178.640 166.380 179.760 ;
  LAYER metal2 ;
  RECT 162.840 178.640 166.380 179.760 ;
  LAYER metal1 ;
  RECT 162.840 178.640 166.380 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 149.200 178.640 152.740 179.760 ;
  LAYER metal4 ;
  RECT 149.200 178.640 152.740 179.760 ;
  LAYER metal3 ;
  RECT 149.200 178.640 152.740 179.760 ;
  LAYER metal2 ;
  RECT 149.200 178.640 152.740 179.760 ;
  LAYER metal1 ;
  RECT 149.200 178.640 152.740 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 82.240 178.640 85.780 179.760 ;
  LAYER metal4 ;
  RECT 82.240 178.640 85.780 179.760 ;
  LAYER metal3 ;
  RECT 82.240 178.640 85.780 179.760 ;
  LAYER metal2 ;
  RECT 82.240 178.640 85.780 179.760 ;
  LAYER metal1 ;
  RECT 82.240 178.640 85.780 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 68.600 178.640 72.140 179.760 ;
  LAYER metal4 ;
  RECT 68.600 178.640 72.140 179.760 ;
  LAYER metal3 ;
  RECT 68.600 178.640 72.140 179.760 ;
  LAYER metal2 ;
  RECT 68.600 178.640 72.140 179.760 ;
  LAYER metal1 ;
  RECT 68.600 178.640 72.140 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 54.960 178.640 58.500 179.760 ;
  LAYER metal4 ;
  RECT 54.960 178.640 58.500 179.760 ;
  LAYER metal3 ;
  RECT 54.960 178.640 58.500 179.760 ;
  LAYER metal2 ;
  RECT 54.960 178.640 58.500 179.760 ;
  LAYER metal1 ;
  RECT 54.960 178.640 58.500 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 41.940 178.640 45.480 179.760 ;
  LAYER metal4 ;
  RECT 41.940 178.640 45.480 179.760 ;
  LAYER metal3 ;
  RECT 41.940 178.640 45.480 179.760 ;
  LAYER metal2 ;
  RECT 41.940 178.640 45.480 179.760 ;
  LAYER metal1 ;
  RECT 41.940 178.640 45.480 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 28.300 178.640 31.840 179.760 ;
  LAYER metal4 ;
  RECT 28.300 178.640 31.840 179.760 ;
  LAYER metal3 ;
  RECT 28.300 178.640 31.840 179.760 ;
  LAYER metal2 ;
  RECT 28.300 178.640 31.840 179.760 ;
  LAYER metal1 ;
  RECT 28.300 178.640 31.840 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 17.140 178.640 20.680 179.760 ;
  LAYER metal4 ;
  RECT 17.140 178.640 20.680 179.760 ;
  LAYER metal3 ;
  RECT 17.140 178.640 20.680 179.760 ;
  LAYER metal2 ;
  RECT 17.140 178.640 20.680 179.760 ;
  LAYER metal1 ;
  RECT 17.140 178.640 20.680 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3531.300 0.000 3534.840 1.120 ;
  LAYER metal4 ;
  RECT 3531.300 0.000 3534.840 1.120 ;
  LAYER metal3 ;
  RECT 3531.300 0.000 3534.840 1.120 ;
  LAYER metal2 ;
  RECT 3531.300 0.000 3534.840 1.120 ;
  LAYER metal1 ;
  RECT 3531.300 0.000 3534.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3517.660 0.000 3521.200 1.120 ;
  LAYER metal4 ;
  RECT 3517.660 0.000 3521.200 1.120 ;
  LAYER metal3 ;
  RECT 3517.660 0.000 3521.200 1.120 ;
  LAYER metal2 ;
  RECT 3517.660 0.000 3521.200 1.120 ;
  LAYER metal1 ;
  RECT 3517.660 0.000 3521.200 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3450.700 0.000 3454.240 1.120 ;
  LAYER metal4 ;
  RECT 3450.700 0.000 3454.240 1.120 ;
  LAYER metal3 ;
  RECT 3450.700 0.000 3454.240 1.120 ;
  LAYER metal2 ;
  RECT 3450.700 0.000 3454.240 1.120 ;
  LAYER metal1 ;
  RECT 3450.700 0.000 3454.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3437.060 0.000 3440.600 1.120 ;
  LAYER metal4 ;
  RECT 3437.060 0.000 3440.600 1.120 ;
  LAYER metal3 ;
  RECT 3437.060 0.000 3440.600 1.120 ;
  LAYER metal2 ;
  RECT 3437.060 0.000 3440.600 1.120 ;
  LAYER metal1 ;
  RECT 3437.060 0.000 3440.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3423.420 0.000 3426.960 1.120 ;
  LAYER metal4 ;
  RECT 3423.420 0.000 3426.960 1.120 ;
  LAYER metal3 ;
  RECT 3423.420 0.000 3426.960 1.120 ;
  LAYER metal2 ;
  RECT 3423.420 0.000 3426.960 1.120 ;
  LAYER metal1 ;
  RECT 3423.420 0.000 3426.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3410.400 0.000 3413.940 1.120 ;
  LAYER metal4 ;
  RECT 3410.400 0.000 3413.940 1.120 ;
  LAYER metal3 ;
  RECT 3410.400 0.000 3413.940 1.120 ;
  LAYER metal2 ;
  RECT 3410.400 0.000 3413.940 1.120 ;
  LAYER metal1 ;
  RECT 3410.400 0.000 3413.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3396.760 0.000 3400.300 1.120 ;
  LAYER metal4 ;
  RECT 3396.760 0.000 3400.300 1.120 ;
  LAYER metal3 ;
  RECT 3396.760 0.000 3400.300 1.120 ;
  LAYER metal2 ;
  RECT 3396.760 0.000 3400.300 1.120 ;
  LAYER metal1 ;
  RECT 3396.760 0.000 3400.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3383.120 0.000 3386.660 1.120 ;
  LAYER metal4 ;
  RECT 3383.120 0.000 3386.660 1.120 ;
  LAYER metal3 ;
  RECT 3383.120 0.000 3386.660 1.120 ;
  LAYER metal2 ;
  RECT 3383.120 0.000 3386.660 1.120 ;
  LAYER metal1 ;
  RECT 3383.120 0.000 3386.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3316.160 0.000 3319.700 1.120 ;
  LAYER metal4 ;
  RECT 3316.160 0.000 3319.700 1.120 ;
  LAYER metal3 ;
  RECT 3316.160 0.000 3319.700 1.120 ;
  LAYER metal2 ;
  RECT 3316.160 0.000 3319.700 1.120 ;
  LAYER metal1 ;
  RECT 3316.160 0.000 3319.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3302.520 0.000 3306.060 1.120 ;
  LAYER metal4 ;
  RECT 3302.520 0.000 3306.060 1.120 ;
  LAYER metal3 ;
  RECT 3302.520 0.000 3306.060 1.120 ;
  LAYER metal2 ;
  RECT 3302.520 0.000 3306.060 1.120 ;
  LAYER metal1 ;
  RECT 3302.520 0.000 3306.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3288.880 0.000 3292.420 1.120 ;
  LAYER metal4 ;
  RECT 3288.880 0.000 3292.420 1.120 ;
  LAYER metal3 ;
  RECT 3288.880 0.000 3292.420 1.120 ;
  LAYER metal2 ;
  RECT 3288.880 0.000 3292.420 1.120 ;
  LAYER metal1 ;
  RECT 3288.880 0.000 3292.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3275.860 0.000 3279.400 1.120 ;
  LAYER metal4 ;
  RECT 3275.860 0.000 3279.400 1.120 ;
  LAYER metal3 ;
  RECT 3275.860 0.000 3279.400 1.120 ;
  LAYER metal2 ;
  RECT 3275.860 0.000 3279.400 1.120 ;
  LAYER metal1 ;
  RECT 3275.860 0.000 3279.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3262.220 0.000 3265.760 1.120 ;
  LAYER metal4 ;
  RECT 3262.220 0.000 3265.760 1.120 ;
  LAYER metal3 ;
  RECT 3262.220 0.000 3265.760 1.120 ;
  LAYER metal2 ;
  RECT 3262.220 0.000 3265.760 1.120 ;
  LAYER metal1 ;
  RECT 3262.220 0.000 3265.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3248.580 0.000 3252.120 1.120 ;
  LAYER metal4 ;
  RECT 3248.580 0.000 3252.120 1.120 ;
  LAYER metal3 ;
  RECT 3248.580 0.000 3252.120 1.120 ;
  LAYER metal2 ;
  RECT 3248.580 0.000 3252.120 1.120 ;
  LAYER metal1 ;
  RECT 3248.580 0.000 3252.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3181.620 0.000 3185.160 1.120 ;
  LAYER metal4 ;
  RECT 3181.620 0.000 3185.160 1.120 ;
  LAYER metal3 ;
  RECT 3181.620 0.000 3185.160 1.120 ;
  LAYER metal2 ;
  RECT 3181.620 0.000 3185.160 1.120 ;
  LAYER metal1 ;
  RECT 3181.620 0.000 3185.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3167.980 0.000 3171.520 1.120 ;
  LAYER metal4 ;
  RECT 3167.980 0.000 3171.520 1.120 ;
  LAYER metal3 ;
  RECT 3167.980 0.000 3171.520 1.120 ;
  LAYER metal2 ;
  RECT 3167.980 0.000 3171.520 1.120 ;
  LAYER metal1 ;
  RECT 3167.980 0.000 3171.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3154.960 0.000 3158.500 1.120 ;
  LAYER metal4 ;
  RECT 3154.960 0.000 3158.500 1.120 ;
  LAYER metal3 ;
  RECT 3154.960 0.000 3158.500 1.120 ;
  LAYER metal2 ;
  RECT 3154.960 0.000 3158.500 1.120 ;
  LAYER metal1 ;
  RECT 3154.960 0.000 3158.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3141.320 0.000 3144.860 1.120 ;
  LAYER metal4 ;
  RECT 3141.320 0.000 3144.860 1.120 ;
  LAYER metal3 ;
  RECT 3141.320 0.000 3144.860 1.120 ;
  LAYER metal2 ;
  RECT 3141.320 0.000 3144.860 1.120 ;
  LAYER metal1 ;
  RECT 3141.320 0.000 3144.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3127.680 0.000 3131.220 1.120 ;
  LAYER metal4 ;
  RECT 3127.680 0.000 3131.220 1.120 ;
  LAYER metal3 ;
  RECT 3127.680 0.000 3131.220 1.120 ;
  LAYER metal2 ;
  RECT 3127.680 0.000 3131.220 1.120 ;
  LAYER metal1 ;
  RECT 3127.680 0.000 3131.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3116.520 0.000 3120.060 1.120 ;
  LAYER metal4 ;
  RECT 3116.520 0.000 3120.060 1.120 ;
  LAYER metal3 ;
  RECT 3116.520 0.000 3120.060 1.120 ;
  LAYER metal2 ;
  RECT 3116.520 0.000 3120.060 1.120 ;
  LAYER metal1 ;
  RECT 3116.520 0.000 3120.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3047.080 0.000 3050.620 1.120 ;
  LAYER metal4 ;
  RECT 3047.080 0.000 3050.620 1.120 ;
  LAYER metal3 ;
  RECT 3047.080 0.000 3050.620 1.120 ;
  LAYER metal2 ;
  RECT 3047.080 0.000 3050.620 1.120 ;
  LAYER metal1 ;
  RECT 3047.080 0.000 3050.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3034.060 0.000 3037.600 1.120 ;
  LAYER metal4 ;
  RECT 3034.060 0.000 3037.600 1.120 ;
  LAYER metal3 ;
  RECT 3034.060 0.000 3037.600 1.120 ;
  LAYER metal2 ;
  RECT 3034.060 0.000 3037.600 1.120 ;
  LAYER metal1 ;
  RECT 3034.060 0.000 3037.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3020.420 0.000 3023.960 1.120 ;
  LAYER metal4 ;
  RECT 3020.420 0.000 3023.960 1.120 ;
  LAYER metal3 ;
  RECT 3020.420 0.000 3023.960 1.120 ;
  LAYER metal2 ;
  RECT 3020.420 0.000 3023.960 1.120 ;
  LAYER metal1 ;
  RECT 3020.420 0.000 3023.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3006.780 0.000 3010.320 1.120 ;
  LAYER metal4 ;
  RECT 3006.780 0.000 3010.320 1.120 ;
  LAYER metal3 ;
  RECT 3006.780 0.000 3010.320 1.120 ;
  LAYER metal2 ;
  RECT 3006.780 0.000 3010.320 1.120 ;
  LAYER metal1 ;
  RECT 3006.780 0.000 3010.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2993.760 0.000 2997.300 1.120 ;
  LAYER metal4 ;
  RECT 2993.760 0.000 2997.300 1.120 ;
  LAYER metal3 ;
  RECT 2993.760 0.000 2997.300 1.120 ;
  LAYER metal2 ;
  RECT 2993.760 0.000 2997.300 1.120 ;
  LAYER metal1 ;
  RECT 2993.760 0.000 2997.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2980.120 0.000 2983.660 1.120 ;
  LAYER metal4 ;
  RECT 2980.120 0.000 2983.660 1.120 ;
  LAYER metal3 ;
  RECT 2980.120 0.000 2983.660 1.120 ;
  LAYER metal2 ;
  RECT 2980.120 0.000 2983.660 1.120 ;
  LAYER metal1 ;
  RECT 2980.120 0.000 2983.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2912.540 0.000 2916.080 1.120 ;
  LAYER metal4 ;
  RECT 2912.540 0.000 2916.080 1.120 ;
  LAYER metal3 ;
  RECT 2912.540 0.000 2916.080 1.120 ;
  LAYER metal2 ;
  RECT 2912.540 0.000 2916.080 1.120 ;
  LAYER metal1 ;
  RECT 2912.540 0.000 2916.080 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2899.520 0.000 2903.060 1.120 ;
  LAYER metal4 ;
  RECT 2899.520 0.000 2903.060 1.120 ;
  LAYER metal3 ;
  RECT 2899.520 0.000 2903.060 1.120 ;
  LAYER metal2 ;
  RECT 2899.520 0.000 2903.060 1.120 ;
  LAYER metal1 ;
  RECT 2899.520 0.000 2903.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2885.880 0.000 2889.420 1.120 ;
  LAYER metal4 ;
  RECT 2885.880 0.000 2889.420 1.120 ;
  LAYER metal3 ;
  RECT 2885.880 0.000 2889.420 1.120 ;
  LAYER metal2 ;
  RECT 2885.880 0.000 2889.420 1.120 ;
  LAYER metal1 ;
  RECT 2885.880 0.000 2889.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2872.240 0.000 2875.780 1.120 ;
  LAYER metal4 ;
  RECT 2872.240 0.000 2875.780 1.120 ;
  LAYER metal3 ;
  RECT 2872.240 0.000 2875.780 1.120 ;
  LAYER metal2 ;
  RECT 2872.240 0.000 2875.780 1.120 ;
  LAYER metal1 ;
  RECT 2872.240 0.000 2875.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2859.220 0.000 2862.760 1.120 ;
  LAYER metal4 ;
  RECT 2859.220 0.000 2862.760 1.120 ;
  LAYER metal3 ;
  RECT 2859.220 0.000 2862.760 1.120 ;
  LAYER metal2 ;
  RECT 2859.220 0.000 2862.760 1.120 ;
  LAYER metal1 ;
  RECT 2859.220 0.000 2862.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2845.580 0.000 2849.120 1.120 ;
  LAYER metal4 ;
  RECT 2845.580 0.000 2849.120 1.120 ;
  LAYER metal3 ;
  RECT 2845.580 0.000 2849.120 1.120 ;
  LAYER metal2 ;
  RECT 2845.580 0.000 2849.120 1.120 ;
  LAYER metal1 ;
  RECT 2845.580 0.000 2849.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2778.620 0.000 2782.160 1.120 ;
  LAYER metal4 ;
  RECT 2778.620 0.000 2782.160 1.120 ;
  LAYER metal3 ;
  RECT 2778.620 0.000 2782.160 1.120 ;
  LAYER metal2 ;
  RECT 2778.620 0.000 2782.160 1.120 ;
  LAYER metal1 ;
  RECT 2778.620 0.000 2782.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2764.980 0.000 2768.520 1.120 ;
  LAYER metal4 ;
  RECT 2764.980 0.000 2768.520 1.120 ;
  LAYER metal3 ;
  RECT 2764.980 0.000 2768.520 1.120 ;
  LAYER metal2 ;
  RECT 2764.980 0.000 2768.520 1.120 ;
  LAYER metal1 ;
  RECT 2764.980 0.000 2768.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2751.340 0.000 2754.880 1.120 ;
  LAYER metal4 ;
  RECT 2751.340 0.000 2754.880 1.120 ;
  LAYER metal3 ;
  RECT 2751.340 0.000 2754.880 1.120 ;
  LAYER metal2 ;
  RECT 2751.340 0.000 2754.880 1.120 ;
  LAYER metal1 ;
  RECT 2751.340 0.000 2754.880 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2738.320 0.000 2741.860 1.120 ;
  LAYER metal4 ;
  RECT 2738.320 0.000 2741.860 1.120 ;
  LAYER metal3 ;
  RECT 2738.320 0.000 2741.860 1.120 ;
  LAYER metal2 ;
  RECT 2738.320 0.000 2741.860 1.120 ;
  LAYER metal1 ;
  RECT 2738.320 0.000 2741.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2724.680 0.000 2728.220 1.120 ;
  LAYER metal4 ;
  RECT 2724.680 0.000 2728.220 1.120 ;
  LAYER metal3 ;
  RECT 2724.680 0.000 2728.220 1.120 ;
  LAYER metal2 ;
  RECT 2724.680 0.000 2728.220 1.120 ;
  LAYER metal1 ;
  RECT 2724.680 0.000 2728.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2711.040 0.000 2714.580 1.120 ;
  LAYER metal4 ;
  RECT 2711.040 0.000 2714.580 1.120 ;
  LAYER metal3 ;
  RECT 2711.040 0.000 2714.580 1.120 ;
  LAYER metal2 ;
  RECT 2711.040 0.000 2714.580 1.120 ;
  LAYER metal1 ;
  RECT 2711.040 0.000 2714.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2644.080 0.000 2647.620 1.120 ;
  LAYER metal4 ;
  RECT 2644.080 0.000 2647.620 1.120 ;
  LAYER metal3 ;
  RECT 2644.080 0.000 2647.620 1.120 ;
  LAYER metal2 ;
  RECT 2644.080 0.000 2647.620 1.120 ;
  LAYER metal1 ;
  RECT 2644.080 0.000 2647.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2630.440 0.000 2633.980 1.120 ;
  LAYER metal4 ;
  RECT 2630.440 0.000 2633.980 1.120 ;
  LAYER metal3 ;
  RECT 2630.440 0.000 2633.980 1.120 ;
  LAYER metal2 ;
  RECT 2630.440 0.000 2633.980 1.120 ;
  LAYER metal1 ;
  RECT 2630.440 0.000 2633.980 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2617.420 0.000 2620.960 1.120 ;
  LAYER metal4 ;
  RECT 2617.420 0.000 2620.960 1.120 ;
  LAYER metal3 ;
  RECT 2617.420 0.000 2620.960 1.120 ;
  LAYER metal2 ;
  RECT 2617.420 0.000 2620.960 1.120 ;
  LAYER metal1 ;
  RECT 2617.420 0.000 2620.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2603.780 0.000 2607.320 1.120 ;
  LAYER metal4 ;
  RECT 2603.780 0.000 2607.320 1.120 ;
  LAYER metal3 ;
  RECT 2603.780 0.000 2607.320 1.120 ;
  LAYER metal2 ;
  RECT 2603.780 0.000 2607.320 1.120 ;
  LAYER metal1 ;
  RECT 2603.780 0.000 2607.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2590.140 0.000 2593.680 1.120 ;
  LAYER metal4 ;
  RECT 2590.140 0.000 2593.680 1.120 ;
  LAYER metal3 ;
  RECT 2590.140 0.000 2593.680 1.120 ;
  LAYER metal2 ;
  RECT 2590.140 0.000 2593.680 1.120 ;
  LAYER metal1 ;
  RECT 2590.140 0.000 2593.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2577.120 0.000 2580.660 1.120 ;
  LAYER metal4 ;
  RECT 2577.120 0.000 2580.660 1.120 ;
  LAYER metal3 ;
  RECT 2577.120 0.000 2580.660 1.120 ;
  LAYER metal2 ;
  RECT 2577.120 0.000 2580.660 1.120 ;
  LAYER metal1 ;
  RECT 2577.120 0.000 2580.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2509.540 0.000 2513.080 1.120 ;
  LAYER metal4 ;
  RECT 2509.540 0.000 2513.080 1.120 ;
  LAYER metal3 ;
  RECT 2509.540 0.000 2513.080 1.120 ;
  LAYER metal2 ;
  RECT 2509.540 0.000 2513.080 1.120 ;
  LAYER metal1 ;
  RECT 2509.540 0.000 2513.080 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2495.900 0.000 2499.440 1.120 ;
  LAYER metal4 ;
  RECT 2495.900 0.000 2499.440 1.120 ;
  LAYER metal3 ;
  RECT 2495.900 0.000 2499.440 1.120 ;
  LAYER metal2 ;
  RECT 2495.900 0.000 2499.440 1.120 ;
  LAYER metal1 ;
  RECT 2495.900 0.000 2499.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2482.880 0.000 2486.420 1.120 ;
  LAYER metal4 ;
  RECT 2482.880 0.000 2486.420 1.120 ;
  LAYER metal3 ;
  RECT 2482.880 0.000 2486.420 1.120 ;
  LAYER metal2 ;
  RECT 2482.880 0.000 2486.420 1.120 ;
  LAYER metal1 ;
  RECT 2482.880 0.000 2486.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2469.240 0.000 2472.780 1.120 ;
  LAYER metal4 ;
  RECT 2469.240 0.000 2472.780 1.120 ;
  LAYER metal3 ;
  RECT 2469.240 0.000 2472.780 1.120 ;
  LAYER metal2 ;
  RECT 2469.240 0.000 2472.780 1.120 ;
  LAYER metal1 ;
  RECT 2469.240 0.000 2472.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2455.600 0.000 2459.140 1.120 ;
  LAYER metal4 ;
  RECT 2455.600 0.000 2459.140 1.120 ;
  LAYER metal3 ;
  RECT 2455.600 0.000 2459.140 1.120 ;
  LAYER metal2 ;
  RECT 2455.600 0.000 2459.140 1.120 ;
  LAYER metal1 ;
  RECT 2455.600 0.000 2459.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2442.580 0.000 2446.120 1.120 ;
  LAYER metal4 ;
  RECT 2442.580 0.000 2446.120 1.120 ;
  LAYER metal3 ;
  RECT 2442.580 0.000 2446.120 1.120 ;
  LAYER metal2 ;
  RECT 2442.580 0.000 2446.120 1.120 ;
  LAYER metal1 ;
  RECT 2442.580 0.000 2446.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2375.000 0.000 2378.540 1.120 ;
  LAYER metal4 ;
  RECT 2375.000 0.000 2378.540 1.120 ;
  LAYER metal3 ;
  RECT 2375.000 0.000 2378.540 1.120 ;
  LAYER metal2 ;
  RECT 2375.000 0.000 2378.540 1.120 ;
  LAYER metal1 ;
  RECT 2375.000 0.000 2378.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2361.980 0.000 2365.520 1.120 ;
  LAYER metal4 ;
  RECT 2361.980 0.000 2365.520 1.120 ;
  LAYER metal3 ;
  RECT 2361.980 0.000 2365.520 1.120 ;
  LAYER metal2 ;
  RECT 2361.980 0.000 2365.520 1.120 ;
  LAYER metal1 ;
  RECT 2361.980 0.000 2365.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2348.340 0.000 2351.880 1.120 ;
  LAYER metal4 ;
  RECT 2348.340 0.000 2351.880 1.120 ;
  LAYER metal3 ;
  RECT 2348.340 0.000 2351.880 1.120 ;
  LAYER metal2 ;
  RECT 2348.340 0.000 2351.880 1.120 ;
  LAYER metal1 ;
  RECT 2348.340 0.000 2351.880 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2334.700 0.000 2338.240 1.120 ;
  LAYER metal4 ;
  RECT 2334.700 0.000 2338.240 1.120 ;
  LAYER metal3 ;
  RECT 2334.700 0.000 2338.240 1.120 ;
  LAYER metal2 ;
  RECT 2334.700 0.000 2338.240 1.120 ;
  LAYER metal1 ;
  RECT 2334.700 0.000 2338.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2321.680 0.000 2325.220 1.120 ;
  LAYER metal4 ;
  RECT 2321.680 0.000 2325.220 1.120 ;
  LAYER metal3 ;
  RECT 2321.680 0.000 2325.220 1.120 ;
  LAYER metal2 ;
  RECT 2321.680 0.000 2325.220 1.120 ;
  LAYER metal1 ;
  RECT 2321.680 0.000 2325.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2308.040 0.000 2311.580 1.120 ;
  LAYER metal4 ;
  RECT 2308.040 0.000 2311.580 1.120 ;
  LAYER metal3 ;
  RECT 2308.040 0.000 2311.580 1.120 ;
  LAYER metal2 ;
  RECT 2308.040 0.000 2311.580 1.120 ;
  LAYER metal1 ;
  RECT 2308.040 0.000 2311.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2241.080 0.000 2244.620 1.120 ;
  LAYER metal4 ;
  RECT 2241.080 0.000 2244.620 1.120 ;
  LAYER metal3 ;
  RECT 2241.080 0.000 2244.620 1.120 ;
  LAYER metal2 ;
  RECT 2241.080 0.000 2244.620 1.120 ;
  LAYER metal1 ;
  RECT 2241.080 0.000 2244.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2227.440 0.000 2230.980 1.120 ;
  LAYER metal4 ;
  RECT 2227.440 0.000 2230.980 1.120 ;
  LAYER metal3 ;
  RECT 2227.440 0.000 2230.980 1.120 ;
  LAYER metal2 ;
  RECT 2227.440 0.000 2230.980 1.120 ;
  LAYER metal1 ;
  RECT 2227.440 0.000 2230.980 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2213.800 0.000 2217.340 1.120 ;
  LAYER metal4 ;
  RECT 2213.800 0.000 2217.340 1.120 ;
  LAYER metal3 ;
  RECT 2213.800 0.000 2217.340 1.120 ;
  LAYER metal2 ;
  RECT 2213.800 0.000 2217.340 1.120 ;
  LAYER metal1 ;
  RECT 2213.800 0.000 2217.340 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2200.780 0.000 2204.320 1.120 ;
  LAYER metal4 ;
  RECT 2200.780 0.000 2204.320 1.120 ;
  LAYER metal3 ;
  RECT 2200.780 0.000 2204.320 1.120 ;
  LAYER metal2 ;
  RECT 2200.780 0.000 2204.320 1.120 ;
  LAYER metal1 ;
  RECT 2200.780 0.000 2204.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2187.140 0.000 2190.680 1.120 ;
  LAYER metal4 ;
  RECT 2187.140 0.000 2190.680 1.120 ;
  LAYER metal3 ;
  RECT 2187.140 0.000 2190.680 1.120 ;
  LAYER metal2 ;
  RECT 2187.140 0.000 2190.680 1.120 ;
  LAYER metal1 ;
  RECT 2187.140 0.000 2190.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2173.500 0.000 2177.040 1.120 ;
  LAYER metal4 ;
  RECT 2173.500 0.000 2177.040 1.120 ;
  LAYER metal3 ;
  RECT 2173.500 0.000 2177.040 1.120 ;
  LAYER metal2 ;
  RECT 2173.500 0.000 2177.040 1.120 ;
  LAYER metal1 ;
  RECT 2173.500 0.000 2177.040 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2106.540 0.000 2110.080 1.120 ;
  LAYER metal4 ;
  RECT 2106.540 0.000 2110.080 1.120 ;
  LAYER metal3 ;
  RECT 2106.540 0.000 2110.080 1.120 ;
  LAYER metal2 ;
  RECT 2106.540 0.000 2110.080 1.120 ;
  LAYER metal1 ;
  RECT 2106.540 0.000 2110.080 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2092.900 0.000 2096.440 1.120 ;
  LAYER metal4 ;
  RECT 2092.900 0.000 2096.440 1.120 ;
  LAYER metal3 ;
  RECT 2092.900 0.000 2096.440 1.120 ;
  LAYER metal2 ;
  RECT 2092.900 0.000 2096.440 1.120 ;
  LAYER metal1 ;
  RECT 2092.900 0.000 2096.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2079.260 0.000 2082.800 1.120 ;
  LAYER metal4 ;
  RECT 2079.260 0.000 2082.800 1.120 ;
  LAYER metal3 ;
  RECT 2079.260 0.000 2082.800 1.120 ;
  LAYER metal2 ;
  RECT 2079.260 0.000 2082.800 1.120 ;
  LAYER metal1 ;
  RECT 2079.260 0.000 2082.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2066.240 0.000 2069.780 1.120 ;
  LAYER metal4 ;
  RECT 2066.240 0.000 2069.780 1.120 ;
  LAYER metal3 ;
  RECT 2066.240 0.000 2069.780 1.120 ;
  LAYER metal2 ;
  RECT 2066.240 0.000 2069.780 1.120 ;
  LAYER metal1 ;
  RECT 2066.240 0.000 2069.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2052.600 0.000 2056.140 1.120 ;
  LAYER metal4 ;
  RECT 2052.600 0.000 2056.140 1.120 ;
  LAYER metal3 ;
  RECT 2052.600 0.000 2056.140 1.120 ;
  LAYER metal2 ;
  RECT 2052.600 0.000 2056.140 1.120 ;
  LAYER metal1 ;
  RECT 2052.600 0.000 2056.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2038.960 0.000 2042.500 1.120 ;
  LAYER metal4 ;
  RECT 2038.960 0.000 2042.500 1.120 ;
  LAYER metal3 ;
  RECT 2038.960 0.000 2042.500 1.120 ;
  LAYER metal2 ;
  RECT 2038.960 0.000 2042.500 1.120 ;
  LAYER metal1 ;
  RECT 2038.960 0.000 2042.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1972.000 0.000 1975.540 1.120 ;
  LAYER metal4 ;
  RECT 1972.000 0.000 1975.540 1.120 ;
  LAYER metal3 ;
  RECT 1972.000 0.000 1975.540 1.120 ;
  LAYER metal2 ;
  RECT 1972.000 0.000 1975.540 1.120 ;
  LAYER metal1 ;
  RECT 1972.000 0.000 1975.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1958.360 0.000 1961.900 1.120 ;
  LAYER metal4 ;
  RECT 1958.360 0.000 1961.900 1.120 ;
  LAYER metal3 ;
  RECT 1958.360 0.000 1961.900 1.120 ;
  LAYER metal2 ;
  RECT 1958.360 0.000 1961.900 1.120 ;
  LAYER metal1 ;
  RECT 1958.360 0.000 1961.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1945.340 0.000 1948.880 1.120 ;
  LAYER metal4 ;
  RECT 1945.340 0.000 1948.880 1.120 ;
  LAYER metal3 ;
  RECT 1945.340 0.000 1948.880 1.120 ;
  LAYER metal2 ;
  RECT 1945.340 0.000 1948.880 1.120 ;
  LAYER metal1 ;
  RECT 1945.340 0.000 1948.880 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1931.700 0.000 1935.240 1.120 ;
  LAYER metal4 ;
  RECT 1931.700 0.000 1935.240 1.120 ;
  LAYER metal3 ;
  RECT 1931.700 0.000 1935.240 1.120 ;
  LAYER metal2 ;
  RECT 1931.700 0.000 1935.240 1.120 ;
  LAYER metal1 ;
  RECT 1931.700 0.000 1935.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1918.060 0.000 1921.600 1.120 ;
  LAYER metal4 ;
  RECT 1918.060 0.000 1921.600 1.120 ;
  LAYER metal3 ;
  RECT 1918.060 0.000 1921.600 1.120 ;
  LAYER metal2 ;
  RECT 1918.060 0.000 1921.600 1.120 ;
  LAYER metal1 ;
  RECT 1918.060 0.000 1921.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1905.040 0.000 1908.580 1.120 ;
  LAYER metal4 ;
  RECT 1905.040 0.000 1908.580 1.120 ;
  LAYER metal3 ;
  RECT 1905.040 0.000 1908.580 1.120 ;
  LAYER metal2 ;
  RECT 1905.040 0.000 1908.580 1.120 ;
  LAYER metal1 ;
  RECT 1905.040 0.000 1908.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1837.460 0.000 1841.000 1.120 ;
  LAYER metal4 ;
  RECT 1837.460 0.000 1841.000 1.120 ;
  LAYER metal3 ;
  RECT 1837.460 0.000 1841.000 1.120 ;
  LAYER metal2 ;
  RECT 1837.460 0.000 1841.000 1.120 ;
  LAYER metal1 ;
  RECT 1837.460 0.000 1841.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1826.300 0.000 1829.840 1.120 ;
  LAYER metal4 ;
  RECT 1826.300 0.000 1829.840 1.120 ;
  LAYER metal3 ;
  RECT 1826.300 0.000 1829.840 1.120 ;
  LAYER metal2 ;
  RECT 1826.300 0.000 1829.840 1.120 ;
  LAYER metal1 ;
  RECT 1826.300 0.000 1829.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1810.180 0.000 1813.720 1.120 ;
  LAYER metal4 ;
  RECT 1810.180 0.000 1813.720 1.120 ;
  LAYER metal3 ;
  RECT 1810.180 0.000 1813.720 1.120 ;
  LAYER metal2 ;
  RECT 1810.180 0.000 1813.720 1.120 ;
  LAYER metal1 ;
  RECT 1810.180 0.000 1813.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1801.500 0.000 1805.040 1.120 ;
  LAYER metal4 ;
  RECT 1801.500 0.000 1805.040 1.120 ;
  LAYER metal3 ;
  RECT 1801.500 0.000 1805.040 1.120 ;
  LAYER metal2 ;
  RECT 1801.500 0.000 1805.040 1.120 ;
  LAYER metal1 ;
  RECT 1801.500 0.000 1805.040 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1792.820 0.000 1796.360 1.120 ;
  LAYER metal4 ;
  RECT 1792.820 0.000 1796.360 1.120 ;
  LAYER metal3 ;
  RECT 1792.820 0.000 1796.360 1.120 ;
  LAYER metal2 ;
  RECT 1792.820 0.000 1796.360 1.120 ;
  LAYER metal1 ;
  RECT 1792.820 0.000 1796.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1779.800 0.000 1783.340 1.120 ;
  LAYER metal4 ;
  RECT 1779.800 0.000 1783.340 1.120 ;
  LAYER metal3 ;
  RECT 1779.800 0.000 1783.340 1.120 ;
  LAYER metal2 ;
  RECT 1779.800 0.000 1783.340 1.120 ;
  LAYER metal1 ;
  RECT 1779.800 0.000 1783.340 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1694.860 0.000 1698.400 1.120 ;
  LAYER metal4 ;
  RECT 1694.860 0.000 1698.400 1.120 ;
  LAYER metal3 ;
  RECT 1694.860 0.000 1698.400 1.120 ;
  LAYER metal2 ;
  RECT 1694.860 0.000 1698.400 1.120 ;
  LAYER metal1 ;
  RECT 1694.860 0.000 1698.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1681.220 0.000 1684.760 1.120 ;
  LAYER metal4 ;
  RECT 1681.220 0.000 1684.760 1.120 ;
  LAYER metal3 ;
  RECT 1681.220 0.000 1684.760 1.120 ;
  LAYER metal2 ;
  RECT 1681.220 0.000 1684.760 1.120 ;
  LAYER metal1 ;
  RECT 1681.220 0.000 1684.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1668.200 0.000 1671.740 1.120 ;
  LAYER metal4 ;
  RECT 1668.200 0.000 1671.740 1.120 ;
  LAYER metal3 ;
  RECT 1668.200 0.000 1671.740 1.120 ;
  LAYER metal2 ;
  RECT 1668.200 0.000 1671.740 1.120 ;
  LAYER metal1 ;
  RECT 1668.200 0.000 1671.740 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1654.560 0.000 1658.100 1.120 ;
  LAYER metal4 ;
  RECT 1654.560 0.000 1658.100 1.120 ;
  LAYER metal3 ;
  RECT 1654.560 0.000 1658.100 1.120 ;
  LAYER metal2 ;
  RECT 1654.560 0.000 1658.100 1.120 ;
  LAYER metal1 ;
  RECT 1654.560 0.000 1658.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1640.920 0.000 1644.460 1.120 ;
  LAYER metal4 ;
  RECT 1640.920 0.000 1644.460 1.120 ;
  LAYER metal3 ;
  RECT 1640.920 0.000 1644.460 1.120 ;
  LAYER metal2 ;
  RECT 1640.920 0.000 1644.460 1.120 ;
  LAYER metal1 ;
  RECT 1640.920 0.000 1644.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1627.900 0.000 1631.440 1.120 ;
  LAYER metal4 ;
  RECT 1627.900 0.000 1631.440 1.120 ;
  LAYER metal3 ;
  RECT 1627.900 0.000 1631.440 1.120 ;
  LAYER metal2 ;
  RECT 1627.900 0.000 1631.440 1.120 ;
  LAYER metal1 ;
  RECT 1627.900 0.000 1631.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1560.320 0.000 1563.860 1.120 ;
  LAYER metal4 ;
  RECT 1560.320 0.000 1563.860 1.120 ;
  LAYER metal3 ;
  RECT 1560.320 0.000 1563.860 1.120 ;
  LAYER metal2 ;
  RECT 1560.320 0.000 1563.860 1.120 ;
  LAYER metal1 ;
  RECT 1560.320 0.000 1563.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1547.300 0.000 1550.840 1.120 ;
  LAYER metal4 ;
  RECT 1547.300 0.000 1550.840 1.120 ;
  LAYER metal3 ;
  RECT 1547.300 0.000 1550.840 1.120 ;
  LAYER metal2 ;
  RECT 1547.300 0.000 1550.840 1.120 ;
  LAYER metal1 ;
  RECT 1547.300 0.000 1550.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1533.660 0.000 1537.200 1.120 ;
  LAYER metal4 ;
  RECT 1533.660 0.000 1537.200 1.120 ;
  LAYER metal3 ;
  RECT 1533.660 0.000 1537.200 1.120 ;
  LAYER metal2 ;
  RECT 1533.660 0.000 1537.200 1.120 ;
  LAYER metal1 ;
  RECT 1533.660 0.000 1537.200 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1520.020 0.000 1523.560 1.120 ;
  LAYER metal4 ;
  RECT 1520.020 0.000 1523.560 1.120 ;
  LAYER metal3 ;
  RECT 1520.020 0.000 1523.560 1.120 ;
  LAYER metal2 ;
  RECT 1520.020 0.000 1523.560 1.120 ;
  LAYER metal1 ;
  RECT 1520.020 0.000 1523.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1507.000 0.000 1510.540 1.120 ;
  LAYER metal4 ;
  RECT 1507.000 0.000 1510.540 1.120 ;
  LAYER metal3 ;
  RECT 1507.000 0.000 1510.540 1.120 ;
  LAYER metal2 ;
  RECT 1507.000 0.000 1510.540 1.120 ;
  LAYER metal1 ;
  RECT 1507.000 0.000 1510.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1493.360 0.000 1496.900 1.120 ;
  LAYER metal4 ;
  RECT 1493.360 0.000 1496.900 1.120 ;
  LAYER metal3 ;
  RECT 1493.360 0.000 1496.900 1.120 ;
  LAYER metal2 ;
  RECT 1493.360 0.000 1496.900 1.120 ;
  LAYER metal1 ;
  RECT 1493.360 0.000 1496.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1426.400 0.000 1429.940 1.120 ;
  LAYER metal4 ;
  RECT 1426.400 0.000 1429.940 1.120 ;
  LAYER metal3 ;
  RECT 1426.400 0.000 1429.940 1.120 ;
  LAYER metal2 ;
  RECT 1426.400 0.000 1429.940 1.120 ;
  LAYER metal1 ;
  RECT 1426.400 0.000 1429.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1412.760 0.000 1416.300 1.120 ;
  LAYER metal4 ;
  RECT 1412.760 0.000 1416.300 1.120 ;
  LAYER metal3 ;
  RECT 1412.760 0.000 1416.300 1.120 ;
  LAYER metal2 ;
  RECT 1412.760 0.000 1416.300 1.120 ;
  LAYER metal1 ;
  RECT 1412.760 0.000 1416.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1399.120 0.000 1402.660 1.120 ;
  LAYER metal4 ;
  RECT 1399.120 0.000 1402.660 1.120 ;
  LAYER metal3 ;
  RECT 1399.120 0.000 1402.660 1.120 ;
  LAYER metal2 ;
  RECT 1399.120 0.000 1402.660 1.120 ;
  LAYER metal1 ;
  RECT 1399.120 0.000 1402.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1386.100 0.000 1389.640 1.120 ;
  LAYER metal4 ;
  RECT 1386.100 0.000 1389.640 1.120 ;
  LAYER metal3 ;
  RECT 1386.100 0.000 1389.640 1.120 ;
  LAYER metal2 ;
  RECT 1386.100 0.000 1389.640 1.120 ;
  LAYER metal1 ;
  RECT 1386.100 0.000 1389.640 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1372.460 0.000 1376.000 1.120 ;
  LAYER metal4 ;
  RECT 1372.460 0.000 1376.000 1.120 ;
  LAYER metal3 ;
  RECT 1372.460 0.000 1376.000 1.120 ;
  LAYER metal2 ;
  RECT 1372.460 0.000 1376.000 1.120 ;
  LAYER metal1 ;
  RECT 1372.460 0.000 1376.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1358.820 0.000 1362.360 1.120 ;
  LAYER metal4 ;
  RECT 1358.820 0.000 1362.360 1.120 ;
  LAYER metal3 ;
  RECT 1358.820 0.000 1362.360 1.120 ;
  LAYER metal2 ;
  RECT 1358.820 0.000 1362.360 1.120 ;
  LAYER metal1 ;
  RECT 1358.820 0.000 1362.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1291.860 0.000 1295.400 1.120 ;
  LAYER metal4 ;
  RECT 1291.860 0.000 1295.400 1.120 ;
  LAYER metal3 ;
  RECT 1291.860 0.000 1295.400 1.120 ;
  LAYER metal2 ;
  RECT 1291.860 0.000 1295.400 1.120 ;
  LAYER metal1 ;
  RECT 1291.860 0.000 1295.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1278.220 0.000 1281.760 1.120 ;
  LAYER metal4 ;
  RECT 1278.220 0.000 1281.760 1.120 ;
  LAYER metal3 ;
  RECT 1278.220 0.000 1281.760 1.120 ;
  LAYER metal2 ;
  RECT 1278.220 0.000 1281.760 1.120 ;
  LAYER metal1 ;
  RECT 1278.220 0.000 1281.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1264.580 0.000 1268.120 1.120 ;
  LAYER metal4 ;
  RECT 1264.580 0.000 1268.120 1.120 ;
  LAYER metal3 ;
  RECT 1264.580 0.000 1268.120 1.120 ;
  LAYER metal2 ;
  RECT 1264.580 0.000 1268.120 1.120 ;
  LAYER metal1 ;
  RECT 1264.580 0.000 1268.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1251.560 0.000 1255.100 1.120 ;
  LAYER metal4 ;
  RECT 1251.560 0.000 1255.100 1.120 ;
  LAYER metal3 ;
  RECT 1251.560 0.000 1255.100 1.120 ;
  LAYER metal2 ;
  RECT 1251.560 0.000 1255.100 1.120 ;
  LAYER metal1 ;
  RECT 1251.560 0.000 1255.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1237.920 0.000 1241.460 1.120 ;
  LAYER metal4 ;
  RECT 1237.920 0.000 1241.460 1.120 ;
  LAYER metal3 ;
  RECT 1237.920 0.000 1241.460 1.120 ;
  LAYER metal2 ;
  RECT 1237.920 0.000 1241.460 1.120 ;
  LAYER metal1 ;
  RECT 1237.920 0.000 1241.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1224.280 0.000 1227.820 1.120 ;
  LAYER metal4 ;
  RECT 1224.280 0.000 1227.820 1.120 ;
  LAYER metal3 ;
  RECT 1224.280 0.000 1227.820 1.120 ;
  LAYER metal2 ;
  RECT 1224.280 0.000 1227.820 1.120 ;
  LAYER metal1 ;
  RECT 1224.280 0.000 1227.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1157.320 0.000 1160.860 1.120 ;
  LAYER metal4 ;
  RECT 1157.320 0.000 1160.860 1.120 ;
  LAYER metal3 ;
  RECT 1157.320 0.000 1160.860 1.120 ;
  LAYER metal2 ;
  RECT 1157.320 0.000 1160.860 1.120 ;
  LAYER metal1 ;
  RECT 1157.320 0.000 1160.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1143.680 0.000 1147.220 1.120 ;
  LAYER metal4 ;
  RECT 1143.680 0.000 1147.220 1.120 ;
  LAYER metal3 ;
  RECT 1143.680 0.000 1147.220 1.120 ;
  LAYER metal2 ;
  RECT 1143.680 0.000 1147.220 1.120 ;
  LAYER metal1 ;
  RECT 1143.680 0.000 1147.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1130.660 0.000 1134.200 1.120 ;
  LAYER metal4 ;
  RECT 1130.660 0.000 1134.200 1.120 ;
  LAYER metal3 ;
  RECT 1130.660 0.000 1134.200 1.120 ;
  LAYER metal2 ;
  RECT 1130.660 0.000 1134.200 1.120 ;
  LAYER metal1 ;
  RECT 1130.660 0.000 1134.200 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1117.020 0.000 1120.560 1.120 ;
  LAYER metal4 ;
  RECT 1117.020 0.000 1120.560 1.120 ;
  LAYER metal3 ;
  RECT 1117.020 0.000 1120.560 1.120 ;
  LAYER metal2 ;
  RECT 1117.020 0.000 1120.560 1.120 ;
  LAYER metal1 ;
  RECT 1117.020 0.000 1120.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1103.380 0.000 1106.920 1.120 ;
  LAYER metal4 ;
  RECT 1103.380 0.000 1106.920 1.120 ;
  LAYER metal3 ;
  RECT 1103.380 0.000 1106.920 1.120 ;
  LAYER metal2 ;
  RECT 1103.380 0.000 1106.920 1.120 ;
  LAYER metal1 ;
  RECT 1103.380 0.000 1106.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1090.360 0.000 1093.900 1.120 ;
  LAYER metal4 ;
  RECT 1090.360 0.000 1093.900 1.120 ;
  LAYER metal3 ;
  RECT 1090.360 0.000 1093.900 1.120 ;
  LAYER metal2 ;
  RECT 1090.360 0.000 1093.900 1.120 ;
  LAYER metal1 ;
  RECT 1090.360 0.000 1093.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1022.780 0.000 1026.320 1.120 ;
  LAYER metal4 ;
  RECT 1022.780 0.000 1026.320 1.120 ;
  LAYER metal3 ;
  RECT 1022.780 0.000 1026.320 1.120 ;
  LAYER metal2 ;
  RECT 1022.780 0.000 1026.320 1.120 ;
  LAYER metal1 ;
  RECT 1022.780 0.000 1026.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1009.760 0.000 1013.300 1.120 ;
  LAYER metal4 ;
  RECT 1009.760 0.000 1013.300 1.120 ;
  LAYER metal3 ;
  RECT 1009.760 0.000 1013.300 1.120 ;
  LAYER metal2 ;
  RECT 1009.760 0.000 1013.300 1.120 ;
  LAYER metal1 ;
  RECT 1009.760 0.000 1013.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 996.120 0.000 999.660 1.120 ;
  LAYER metal4 ;
  RECT 996.120 0.000 999.660 1.120 ;
  LAYER metal3 ;
  RECT 996.120 0.000 999.660 1.120 ;
  LAYER metal2 ;
  RECT 996.120 0.000 999.660 1.120 ;
  LAYER metal1 ;
  RECT 996.120 0.000 999.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 982.480 0.000 986.020 1.120 ;
  LAYER metal4 ;
  RECT 982.480 0.000 986.020 1.120 ;
  LAYER metal3 ;
  RECT 982.480 0.000 986.020 1.120 ;
  LAYER metal2 ;
  RECT 982.480 0.000 986.020 1.120 ;
  LAYER metal1 ;
  RECT 982.480 0.000 986.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 969.460 0.000 973.000 1.120 ;
  LAYER metal4 ;
  RECT 969.460 0.000 973.000 1.120 ;
  LAYER metal3 ;
  RECT 969.460 0.000 973.000 1.120 ;
  LAYER metal2 ;
  RECT 969.460 0.000 973.000 1.120 ;
  LAYER metal1 ;
  RECT 969.460 0.000 973.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 955.820 0.000 959.360 1.120 ;
  LAYER metal4 ;
  RECT 955.820 0.000 959.360 1.120 ;
  LAYER metal3 ;
  RECT 955.820 0.000 959.360 1.120 ;
  LAYER metal2 ;
  RECT 955.820 0.000 959.360 1.120 ;
  LAYER metal1 ;
  RECT 955.820 0.000 959.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 888.240 0.000 891.780 1.120 ;
  LAYER metal4 ;
  RECT 888.240 0.000 891.780 1.120 ;
  LAYER metal3 ;
  RECT 888.240 0.000 891.780 1.120 ;
  LAYER metal2 ;
  RECT 888.240 0.000 891.780 1.120 ;
  LAYER metal1 ;
  RECT 888.240 0.000 891.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 877.080 0.000 880.620 1.120 ;
  LAYER metal4 ;
  RECT 877.080 0.000 880.620 1.120 ;
  LAYER metal3 ;
  RECT 877.080 0.000 880.620 1.120 ;
  LAYER metal2 ;
  RECT 877.080 0.000 880.620 1.120 ;
  LAYER metal1 ;
  RECT 877.080 0.000 880.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 861.580 0.000 865.120 1.120 ;
  LAYER metal4 ;
  RECT 861.580 0.000 865.120 1.120 ;
  LAYER metal3 ;
  RECT 861.580 0.000 865.120 1.120 ;
  LAYER metal2 ;
  RECT 861.580 0.000 865.120 1.120 ;
  LAYER metal1 ;
  RECT 861.580 0.000 865.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 847.940 0.000 851.480 1.120 ;
  LAYER metal4 ;
  RECT 847.940 0.000 851.480 1.120 ;
  LAYER metal3 ;
  RECT 847.940 0.000 851.480 1.120 ;
  LAYER metal2 ;
  RECT 847.940 0.000 851.480 1.120 ;
  LAYER metal1 ;
  RECT 847.940 0.000 851.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 834.920 0.000 838.460 1.120 ;
  LAYER metal4 ;
  RECT 834.920 0.000 838.460 1.120 ;
  LAYER metal3 ;
  RECT 834.920 0.000 838.460 1.120 ;
  LAYER metal2 ;
  RECT 834.920 0.000 838.460 1.120 ;
  LAYER metal1 ;
  RECT 834.920 0.000 838.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 821.280 0.000 824.820 1.120 ;
  LAYER metal4 ;
  RECT 821.280 0.000 824.820 1.120 ;
  LAYER metal3 ;
  RECT 821.280 0.000 824.820 1.120 ;
  LAYER metal2 ;
  RECT 821.280 0.000 824.820 1.120 ;
  LAYER metal1 ;
  RECT 821.280 0.000 824.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 754.320 0.000 757.860 1.120 ;
  LAYER metal4 ;
  RECT 754.320 0.000 757.860 1.120 ;
  LAYER metal3 ;
  RECT 754.320 0.000 757.860 1.120 ;
  LAYER metal2 ;
  RECT 754.320 0.000 757.860 1.120 ;
  LAYER metal1 ;
  RECT 754.320 0.000 757.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 740.680 0.000 744.220 1.120 ;
  LAYER metal4 ;
  RECT 740.680 0.000 744.220 1.120 ;
  LAYER metal3 ;
  RECT 740.680 0.000 744.220 1.120 ;
  LAYER metal2 ;
  RECT 740.680 0.000 744.220 1.120 ;
  LAYER metal1 ;
  RECT 740.680 0.000 744.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 727.040 0.000 730.580 1.120 ;
  LAYER metal4 ;
  RECT 727.040 0.000 730.580 1.120 ;
  LAYER metal3 ;
  RECT 727.040 0.000 730.580 1.120 ;
  LAYER metal2 ;
  RECT 727.040 0.000 730.580 1.120 ;
  LAYER metal1 ;
  RECT 727.040 0.000 730.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 714.020 0.000 717.560 1.120 ;
  LAYER metal4 ;
  RECT 714.020 0.000 717.560 1.120 ;
  LAYER metal3 ;
  RECT 714.020 0.000 717.560 1.120 ;
  LAYER metal2 ;
  RECT 714.020 0.000 717.560 1.120 ;
  LAYER metal1 ;
  RECT 714.020 0.000 717.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 700.380 0.000 703.920 1.120 ;
  LAYER metal4 ;
  RECT 700.380 0.000 703.920 1.120 ;
  LAYER metal3 ;
  RECT 700.380 0.000 703.920 1.120 ;
  LAYER metal2 ;
  RECT 700.380 0.000 703.920 1.120 ;
  LAYER metal1 ;
  RECT 700.380 0.000 703.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 686.740 0.000 690.280 1.120 ;
  LAYER metal4 ;
  RECT 686.740 0.000 690.280 1.120 ;
  LAYER metal3 ;
  RECT 686.740 0.000 690.280 1.120 ;
  LAYER metal2 ;
  RECT 686.740 0.000 690.280 1.120 ;
  LAYER metal1 ;
  RECT 686.740 0.000 690.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 619.780 0.000 623.320 1.120 ;
  LAYER metal4 ;
  RECT 619.780 0.000 623.320 1.120 ;
  LAYER metal3 ;
  RECT 619.780 0.000 623.320 1.120 ;
  LAYER metal2 ;
  RECT 619.780 0.000 623.320 1.120 ;
  LAYER metal1 ;
  RECT 619.780 0.000 623.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 606.140 0.000 609.680 1.120 ;
  LAYER metal4 ;
  RECT 606.140 0.000 609.680 1.120 ;
  LAYER metal3 ;
  RECT 606.140 0.000 609.680 1.120 ;
  LAYER metal2 ;
  RECT 606.140 0.000 609.680 1.120 ;
  LAYER metal1 ;
  RECT 606.140 0.000 609.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 593.120 0.000 596.660 1.120 ;
  LAYER metal4 ;
  RECT 593.120 0.000 596.660 1.120 ;
  LAYER metal3 ;
  RECT 593.120 0.000 596.660 1.120 ;
  LAYER metal2 ;
  RECT 593.120 0.000 596.660 1.120 ;
  LAYER metal1 ;
  RECT 593.120 0.000 596.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 579.480 0.000 583.020 1.120 ;
  LAYER metal4 ;
  RECT 579.480 0.000 583.020 1.120 ;
  LAYER metal3 ;
  RECT 579.480 0.000 583.020 1.120 ;
  LAYER metal2 ;
  RECT 579.480 0.000 583.020 1.120 ;
  LAYER metal1 ;
  RECT 579.480 0.000 583.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER metal4 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER metal3 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER metal2 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER metal1 ;
  RECT 565.840 0.000 569.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 552.820 0.000 556.360 1.120 ;
  LAYER metal4 ;
  RECT 552.820 0.000 556.360 1.120 ;
  LAYER metal3 ;
  RECT 552.820 0.000 556.360 1.120 ;
  LAYER metal2 ;
  RECT 552.820 0.000 556.360 1.120 ;
  LAYER metal1 ;
  RECT 552.820 0.000 556.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 485.240 0.000 488.780 1.120 ;
  LAYER metal4 ;
  RECT 485.240 0.000 488.780 1.120 ;
  LAYER metal3 ;
  RECT 485.240 0.000 488.780 1.120 ;
  LAYER metal2 ;
  RECT 485.240 0.000 488.780 1.120 ;
  LAYER metal1 ;
  RECT 485.240 0.000 488.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 471.600 0.000 475.140 1.120 ;
  LAYER metal4 ;
  RECT 471.600 0.000 475.140 1.120 ;
  LAYER metal3 ;
  RECT 471.600 0.000 475.140 1.120 ;
  LAYER metal2 ;
  RECT 471.600 0.000 475.140 1.120 ;
  LAYER metal1 ;
  RECT 471.600 0.000 475.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 458.580 0.000 462.120 1.120 ;
  LAYER metal4 ;
  RECT 458.580 0.000 462.120 1.120 ;
  LAYER metal3 ;
  RECT 458.580 0.000 462.120 1.120 ;
  LAYER metal2 ;
  RECT 458.580 0.000 462.120 1.120 ;
  LAYER metal1 ;
  RECT 458.580 0.000 462.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 447.420 0.000 450.960 1.120 ;
  LAYER metal4 ;
  RECT 447.420 0.000 450.960 1.120 ;
  LAYER metal3 ;
  RECT 447.420 0.000 450.960 1.120 ;
  LAYER metal2 ;
  RECT 447.420 0.000 450.960 1.120 ;
  LAYER metal1 ;
  RECT 447.420 0.000 450.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER metal4 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER metal3 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER metal2 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER metal1 ;
  RECT 431.300 0.000 434.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 418.280 0.000 421.820 1.120 ;
  LAYER metal4 ;
  RECT 418.280 0.000 421.820 1.120 ;
  LAYER metal3 ;
  RECT 418.280 0.000 421.820 1.120 ;
  LAYER metal2 ;
  RECT 418.280 0.000 421.820 1.120 ;
  LAYER metal1 ;
  RECT 418.280 0.000 421.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 350.700 0.000 354.240 1.120 ;
  LAYER metal4 ;
  RECT 350.700 0.000 354.240 1.120 ;
  LAYER metal3 ;
  RECT 350.700 0.000 354.240 1.120 ;
  LAYER metal2 ;
  RECT 350.700 0.000 354.240 1.120 ;
  LAYER metal1 ;
  RECT 350.700 0.000 354.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 337.680 0.000 341.220 1.120 ;
  LAYER metal4 ;
  RECT 337.680 0.000 341.220 1.120 ;
  LAYER metal3 ;
  RECT 337.680 0.000 341.220 1.120 ;
  LAYER metal2 ;
  RECT 337.680 0.000 341.220 1.120 ;
  LAYER metal1 ;
  RECT 337.680 0.000 341.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 324.040 0.000 327.580 1.120 ;
  LAYER metal4 ;
  RECT 324.040 0.000 327.580 1.120 ;
  LAYER metal3 ;
  RECT 324.040 0.000 327.580 1.120 ;
  LAYER metal2 ;
  RECT 324.040 0.000 327.580 1.120 ;
  LAYER metal1 ;
  RECT 324.040 0.000 327.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 310.400 0.000 313.940 1.120 ;
  LAYER metal4 ;
  RECT 310.400 0.000 313.940 1.120 ;
  LAYER metal3 ;
  RECT 310.400 0.000 313.940 1.120 ;
  LAYER metal2 ;
  RECT 310.400 0.000 313.940 1.120 ;
  LAYER metal1 ;
  RECT 310.400 0.000 313.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 297.380 0.000 300.920 1.120 ;
  LAYER metal4 ;
  RECT 297.380 0.000 300.920 1.120 ;
  LAYER metal3 ;
  RECT 297.380 0.000 300.920 1.120 ;
  LAYER metal2 ;
  RECT 297.380 0.000 300.920 1.120 ;
  LAYER metal1 ;
  RECT 297.380 0.000 300.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 283.740 0.000 287.280 1.120 ;
  LAYER metal4 ;
  RECT 283.740 0.000 287.280 1.120 ;
  LAYER metal3 ;
  RECT 283.740 0.000 287.280 1.120 ;
  LAYER metal2 ;
  RECT 283.740 0.000 287.280 1.120 ;
  LAYER metal1 ;
  RECT 283.740 0.000 287.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 216.780 0.000 220.320 1.120 ;
  LAYER metal4 ;
  RECT 216.780 0.000 220.320 1.120 ;
  LAYER metal3 ;
  RECT 216.780 0.000 220.320 1.120 ;
  LAYER metal2 ;
  RECT 216.780 0.000 220.320 1.120 ;
  LAYER metal1 ;
  RECT 216.780 0.000 220.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 203.140 0.000 206.680 1.120 ;
  LAYER metal4 ;
  RECT 203.140 0.000 206.680 1.120 ;
  LAYER metal3 ;
  RECT 203.140 0.000 206.680 1.120 ;
  LAYER metal2 ;
  RECT 203.140 0.000 206.680 1.120 ;
  LAYER metal1 ;
  RECT 203.140 0.000 206.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 189.500 0.000 193.040 1.120 ;
  LAYER metal4 ;
  RECT 189.500 0.000 193.040 1.120 ;
  LAYER metal3 ;
  RECT 189.500 0.000 193.040 1.120 ;
  LAYER metal2 ;
  RECT 189.500 0.000 193.040 1.120 ;
  LAYER metal1 ;
  RECT 189.500 0.000 193.040 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER metal4 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER metal3 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER metal2 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER metal1 ;
  RECT 176.480 0.000 180.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 162.840 0.000 166.380 1.120 ;
  LAYER metal4 ;
  RECT 162.840 0.000 166.380 1.120 ;
  LAYER metal3 ;
  RECT 162.840 0.000 166.380 1.120 ;
  LAYER metal2 ;
  RECT 162.840 0.000 166.380 1.120 ;
  LAYER metal1 ;
  RECT 162.840 0.000 166.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 149.200 0.000 152.740 1.120 ;
  LAYER metal4 ;
  RECT 149.200 0.000 152.740 1.120 ;
  LAYER metal3 ;
  RECT 149.200 0.000 152.740 1.120 ;
  LAYER metal2 ;
  RECT 149.200 0.000 152.740 1.120 ;
  LAYER metal1 ;
  RECT 149.200 0.000 152.740 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 82.240 0.000 85.780 1.120 ;
  LAYER metal4 ;
  RECT 82.240 0.000 85.780 1.120 ;
  LAYER metal3 ;
  RECT 82.240 0.000 85.780 1.120 ;
  LAYER metal2 ;
  RECT 82.240 0.000 85.780 1.120 ;
  LAYER metal1 ;
  RECT 82.240 0.000 85.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 68.600 0.000 72.140 1.120 ;
  LAYER metal4 ;
  RECT 68.600 0.000 72.140 1.120 ;
  LAYER metal3 ;
  RECT 68.600 0.000 72.140 1.120 ;
  LAYER metal2 ;
  RECT 68.600 0.000 72.140 1.120 ;
  LAYER metal1 ;
  RECT 68.600 0.000 72.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER metal4 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER metal3 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER metal2 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER metal1 ;
  RECT 54.960 0.000 58.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER metal4 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER metal3 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER metal2 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER metal1 ;
  RECT 41.940 0.000 45.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER metal4 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER metal3 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER metal2 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER metal1 ;
  RECT 28.300 0.000 31.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 17.140 0.000 20.680 1.120 ;
  LAYER metal4 ;
  RECT 17.140 0.000 20.680 1.120 ;
  LAYER metal3 ;
  RECT 17.140 0.000 20.680 1.120 ;
  LAYER metal2 ;
  RECT 17.140 0.000 20.680 1.120 ;
  LAYER metal1 ;
  RECT 17.140 0.000 20.680 1.120 ;
 END
END GND
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal5 ;
  RECT 3546.520 164.420 3547.640 167.660 ;
  LAYER metal4 ;
  RECT 3546.520 164.420 3547.640 167.660 ;
  LAYER metal3 ;
  RECT 3546.520 164.420 3547.640 167.660 ;
  LAYER metal2 ;
  RECT 3546.520 164.420 3547.640 167.660 ;
  LAYER metal1 ;
  RECT 3546.520 164.420 3547.640 167.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3546.520 125.220 3547.640 128.460 ;
  LAYER metal4 ;
  RECT 3546.520 125.220 3547.640 128.460 ;
  LAYER metal3 ;
  RECT 3546.520 125.220 3547.640 128.460 ;
  LAYER metal2 ;
  RECT 3546.520 125.220 3547.640 128.460 ;
  LAYER metal1 ;
  RECT 3546.520 125.220 3547.640 128.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3546.520 117.380 3547.640 120.620 ;
  LAYER metal4 ;
  RECT 3546.520 117.380 3547.640 120.620 ;
  LAYER metal3 ;
  RECT 3546.520 117.380 3547.640 120.620 ;
  LAYER metal2 ;
  RECT 3546.520 117.380 3547.640 120.620 ;
  LAYER metal1 ;
  RECT 3546.520 117.380 3547.640 120.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3546.520 109.540 3547.640 112.780 ;
  LAYER metal4 ;
  RECT 3546.520 109.540 3547.640 112.780 ;
  LAYER metal3 ;
  RECT 3546.520 109.540 3547.640 112.780 ;
  LAYER metal2 ;
  RECT 3546.520 109.540 3547.640 112.780 ;
  LAYER metal1 ;
  RECT 3546.520 109.540 3547.640 112.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3546.520 101.700 3547.640 104.940 ;
  LAYER metal4 ;
  RECT 3546.520 101.700 3547.640 104.940 ;
  LAYER metal3 ;
  RECT 3546.520 101.700 3547.640 104.940 ;
  LAYER metal2 ;
  RECT 3546.520 101.700 3547.640 104.940 ;
  LAYER metal1 ;
  RECT 3546.520 101.700 3547.640 104.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3546.520 93.860 3547.640 97.100 ;
  LAYER metal4 ;
  RECT 3546.520 93.860 3547.640 97.100 ;
  LAYER metal3 ;
  RECT 3546.520 93.860 3547.640 97.100 ;
  LAYER metal2 ;
  RECT 3546.520 93.860 3547.640 97.100 ;
  LAYER metal1 ;
  RECT 3546.520 93.860 3547.640 97.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3546.520 86.020 3547.640 89.260 ;
  LAYER metal4 ;
  RECT 3546.520 86.020 3547.640 89.260 ;
  LAYER metal3 ;
  RECT 3546.520 86.020 3547.640 89.260 ;
  LAYER metal2 ;
  RECT 3546.520 86.020 3547.640 89.260 ;
  LAYER metal1 ;
  RECT 3546.520 86.020 3547.640 89.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3546.520 46.820 3547.640 50.060 ;
  LAYER metal4 ;
  RECT 3546.520 46.820 3547.640 50.060 ;
  LAYER metal3 ;
  RECT 3546.520 46.820 3547.640 50.060 ;
  LAYER metal2 ;
  RECT 3546.520 46.820 3547.640 50.060 ;
  LAYER metal1 ;
  RECT 3546.520 46.820 3547.640 50.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3546.520 38.980 3547.640 42.220 ;
  LAYER metal4 ;
  RECT 3546.520 38.980 3547.640 42.220 ;
  LAYER metal3 ;
  RECT 3546.520 38.980 3547.640 42.220 ;
  LAYER metal2 ;
  RECT 3546.520 38.980 3547.640 42.220 ;
  LAYER metal1 ;
  RECT 3546.520 38.980 3547.640 42.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3546.520 31.140 3547.640 34.380 ;
  LAYER metal4 ;
  RECT 3546.520 31.140 3547.640 34.380 ;
  LAYER metal3 ;
  RECT 3546.520 31.140 3547.640 34.380 ;
  LAYER metal2 ;
  RECT 3546.520 31.140 3547.640 34.380 ;
  LAYER metal1 ;
  RECT 3546.520 31.140 3547.640 34.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3546.520 23.300 3547.640 26.540 ;
  LAYER metal4 ;
  RECT 3546.520 23.300 3547.640 26.540 ;
  LAYER metal3 ;
  RECT 3546.520 23.300 3547.640 26.540 ;
  LAYER metal2 ;
  RECT 3546.520 23.300 3547.640 26.540 ;
  LAYER metal1 ;
  RECT 3546.520 23.300 3547.640 26.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3546.520 15.460 3547.640 18.700 ;
  LAYER metal4 ;
  RECT 3546.520 15.460 3547.640 18.700 ;
  LAYER metal3 ;
  RECT 3546.520 15.460 3547.640 18.700 ;
  LAYER metal2 ;
  RECT 3546.520 15.460 3547.640 18.700 ;
  LAYER metal1 ;
  RECT 3546.520 15.460 3547.640 18.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3546.520 7.620 3547.640 10.860 ;
  LAYER metal4 ;
  RECT 3546.520 7.620 3547.640 10.860 ;
  LAYER metal3 ;
  RECT 3546.520 7.620 3547.640 10.860 ;
  LAYER metal2 ;
  RECT 3546.520 7.620 3547.640 10.860 ;
  LAYER metal1 ;
  RECT 3546.520 7.620 3547.640 10.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER metal4 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER metal3 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER metal2 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER metal1 ;
  RECT 0.000 164.420 1.120 167.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER metal4 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER metal3 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER metal2 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER metal1 ;
  RECT 0.000 125.220 1.120 128.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER metal4 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER metal3 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER metal2 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER metal1 ;
  RECT 0.000 117.380 1.120 120.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER metal4 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER metal3 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER metal2 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER metal1 ;
  RECT 0.000 109.540 1.120 112.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER metal4 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER metal3 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER metal2 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER metal1 ;
  RECT 0.000 101.700 1.120 104.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER metal4 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER metal3 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER metal2 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER metal1 ;
  RECT 0.000 93.860 1.120 97.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER metal4 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER metal3 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER metal2 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER metal1 ;
  RECT 0.000 86.020 1.120 89.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER metal4 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER metal3 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER metal2 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER metal1 ;
  RECT 0.000 46.820 1.120 50.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER metal4 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER metal3 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER metal2 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER metal1 ;
  RECT 0.000 38.980 1.120 42.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER metal4 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER metal3 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER metal2 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER metal1 ;
  RECT 0.000 31.140 1.120 34.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER metal4 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER metal3 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER metal2 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER metal1 ;
  RECT 0.000 23.300 1.120 26.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER metal4 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER metal3 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER metal2 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER metal1 ;
  RECT 0.000 15.460 1.120 18.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER metal4 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER metal3 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER metal2 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER metal1 ;
  RECT 0.000 7.620 1.120 10.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3535.640 178.640 3539.180 179.760 ;
  LAYER metal4 ;
  RECT 3535.640 178.640 3539.180 179.760 ;
  LAYER metal3 ;
  RECT 3535.640 178.640 3539.180 179.760 ;
  LAYER metal2 ;
  RECT 3535.640 178.640 3539.180 179.760 ;
  LAYER metal1 ;
  RECT 3535.640 178.640 3539.180 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3526.960 178.640 3530.500 179.760 ;
  LAYER metal4 ;
  RECT 3526.960 178.640 3530.500 179.760 ;
  LAYER metal3 ;
  RECT 3526.960 178.640 3530.500 179.760 ;
  LAYER metal2 ;
  RECT 3526.960 178.640 3530.500 179.760 ;
  LAYER metal1 ;
  RECT 3526.960 178.640 3530.500 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3513.320 178.640 3516.860 179.760 ;
  LAYER metal4 ;
  RECT 3513.320 178.640 3516.860 179.760 ;
  LAYER metal3 ;
  RECT 3513.320 178.640 3516.860 179.760 ;
  LAYER metal2 ;
  RECT 3513.320 178.640 3516.860 179.760 ;
  LAYER metal1 ;
  RECT 3513.320 178.640 3516.860 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3446.360 178.640 3449.900 179.760 ;
  LAYER metal4 ;
  RECT 3446.360 178.640 3449.900 179.760 ;
  LAYER metal3 ;
  RECT 3446.360 178.640 3449.900 179.760 ;
  LAYER metal2 ;
  RECT 3446.360 178.640 3449.900 179.760 ;
  LAYER metal1 ;
  RECT 3446.360 178.640 3449.900 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3432.720 178.640 3436.260 179.760 ;
  LAYER metal4 ;
  RECT 3432.720 178.640 3436.260 179.760 ;
  LAYER metal3 ;
  RECT 3432.720 178.640 3436.260 179.760 ;
  LAYER metal2 ;
  RECT 3432.720 178.640 3436.260 179.760 ;
  LAYER metal1 ;
  RECT 3432.720 178.640 3436.260 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3419.080 178.640 3422.620 179.760 ;
  LAYER metal4 ;
  RECT 3419.080 178.640 3422.620 179.760 ;
  LAYER metal3 ;
  RECT 3419.080 178.640 3422.620 179.760 ;
  LAYER metal2 ;
  RECT 3419.080 178.640 3422.620 179.760 ;
  LAYER metal1 ;
  RECT 3419.080 178.640 3422.620 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3406.060 178.640 3409.600 179.760 ;
  LAYER metal4 ;
  RECT 3406.060 178.640 3409.600 179.760 ;
  LAYER metal3 ;
  RECT 3406.060 178.640 3409.600 179.760 ;
  LAYER metal2 ;
  RECT 3406.060 178.640 3409.600 179.760 ;
  LAYER metal1 ;
  RECT 3406.060 178.640 3409.600 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3392.420 178.640 3395.960 179.760 ;
  LAYER metal4 ;
  RECT 3392.420 178.640 3395.960 179.760 ;
  LAYER metal3 ;
  RECT 3392.420 178.640 3395.960 179.760 ;
  LAYER metal2 ;
  RECT 3392.420 178.640 3395.960 179.760 ;
  LAYER metal1 ;
  RECT 3392.420 178.640 3395.960 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3378.780 178.640 3382.320 179.760 ;
  LAYER metal4 ;
  RECT 3378.780 178.640 3382.320 179.760 ;
  LAYER metal3 ;
  RECT 3378.780 178.640 3382.320 179.760 ;
  LAYER metal2 ;
  RECT 3378.780 178.640 3382.320 179.760 ;
  LAYER metal1 ;
  RECT 3378.780 178.640 3382.320 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3311.820 178.640 3315.360 179.760 ;
  LAYER metal4 ;
  RECT 3311.820 178.640 3315.360 179.760 ;
  LAYER metal3 ;
  RECT 3311.820 178.640 3315.360 179.760 ;
  LAYER metal2 ;
  RECT 3311.820 178.640 3315.360 179.760 ;
  LAYER metal1 ;
  RECT 3311.820 178.640 3315.360 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3298.180 178.640 3301.720 179.760 ;
  LAYER metal4 ;
  RECT 3298.180 178.640 3301.720 179.760 ;
  LAYER metal3 ;
  RECT 3298.180 178.640 3301.720 179.760 ;
  LAYER metal2 ;
  RECT 3298.180 178.640 3301.720 179.760 ;
  LAYER metal1 ;
  RECT 3298.180 178.640 3301.720 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3284.540 178.640 3288.080 179.760 ;
  LAYER metal4 ;
  RECT 3284.540 178.640 3288.080 179.760 ;
  LAYER metal3 ;
  RECT 3284.540 178.640 3288.080 179.760 ;
  LAYER metal2 ;
  RECT 3284.540 178.640 3288.080 179.760 ;
  LAYER metal1 ;
  RECT 3284.540 178.640 3288.080 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3271.520 178.640 3275.060 179.760 ;
  LAYER metal4 ;
  RECT 3271.520 178.640 3275.060 179.760 ;
  LAYER metal3 ;
  RECT 3271.520 178.640 3275.060 179.760 ;
  LAYER metal2 ;
  RECT 3271.520 178.640 3275.060 179.760 ;
  LAYER metal1 ;
  RECT 3271.520 178.640 3275.060 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3257.880 178.640 3261.420 179.760 ;
  LAYER metal4 ;
  RECT 3257.880 178.640 3261.420 179.760 ;
  LAYER metal3 ;
  RECT 3257.880 178.640 3261.420 179.760 ;
  LAYER metal2 ;
  RECT 3257.880 178.640 3261.420 179.760 ;
  LAYER metal1 ;
  RECT 3257.880 178.640 3261.420 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3244.240 178.640 3247.780 179.760 ;
  LAYER metal4 ;
  RECT 3244.240 178.640 3247.780 179.760 ;
  LAYER metal3 ;
  RECT 3244.240 178.640 3247.780 179.760 ;
  LAYER metal2 ;
  RECT 3244.240 178.640 3247.780 179.760 ;
  LAYER metal1 ;
  RECT 3244.240 178.640 3247.780 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3177.280 178.640 3180.820 179.760 ;
  LAYER metal4 ;
  RECT 3177.280 178.640 3180.820 179.760 ;
  LAYER metal3 ;
  RECT 3177.280 178.640 3180.820 179.760 ;
  LAYER metal2 ;
  RECT 3177.280 178.640 3180.820 179.760 ;
  LAYER metal1 ;
  RECT 3177.280 178.640 3180.820 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3163.640 178.640 3167.180 179.760 ;
  LAYER metal4 ;
  RECT 3163.640 178.640 3167.180 179.760 ;
  LAYER metal3 ;
  RECT 3163.640 178.640 3167.180 179.760 ;
  LAYER metal2 ;
  RECT 3163.640 178.640 3167.180 179.760 ;
  LAYER metal1 ;
  RECT 3163.640 178.640 3167.180 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3150.620 178.640 3154.160 179.760 ;
  LAYER metal4 ;
  RECT 3150.620 178.640 3154.160 179.760 ;
  LAYER metal3 ;
  RECT 3150.620 178.640 3154.160 179.760 ;
  LAYER metal2 ;
  RECT 3150.620 178.640 3154.160 179.760 ;
  LAYER metal1 ;
  RECT 3150.620 178.640 3154.160 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3136.980 178.640 3140.520 179.760 ;
  LAYER metal4 ;
  RECT 3136.980 178.640 3140.520 179.760 ;
  LAYER metal3 ;
  RECT 3136.980 178.640 3140.520 179.760 ;
  LAYER metal2 ;
  RECT 3136.980 178.640 3140.520 179.760 ;
  LAYER metal1 ;
  RECT 3136.980 178.640 3140.520 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3123.340 178.640 3126.880 179.760 ;
  LAYER metal4 ;
  RECT 3123.340 178.640 3126.880 179.760 ;
  LAYER metal3 ;
  RECT 3123.340 178.640 3126.880 179.760 ;
  LAYER metal2 ;
  RECT 3123.340 178.640 3126.880 179.760 ;
  LAYER metal1 ;
  RECT 3123.340 178.640 3126.880 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3112.180 178.640 3115.720 179.760 ;
  LAYER metal4 ;
  RECT 3112.180 178.640 3115.720 179.760 ;
  LAYER metal3 ;
  RECT 3112.180 178.640 3115.720 179.760 ;
  LAYER metal2 ;
  RECT 3112.180 178.640 3115.720 179.760 ;
  LAYER metal1 ;
  RECT 3112.180 178.640 3115.720 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3042.740 178.640 3046.280 179.760 ;
  LAYER metal4 ;
  RECT 3042.740 178.640 3046.280 179.760 ;
  LAYER metal3 ;
  RECT 3042.740 178.640 3046.280 179.760 ;
  LAYER metal2 ;
  RECT 3042.740 178.640 3046.280 179.760 ;
  LAYER metal1 ;
  RECT 3042.740 178.640 3046.280 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3029.720 178.640 3033.260 179.760 ;
  LAYER metal4 ;
  RECT 3029.720 178.640 3033.260 179.760 ;
  LAYER metal3 ;
  RECT 3029.720 178.640 3033.260 179.760 ;
  LAYER metal2 ;
  RECT 3029.720 178.640 3033.260 179.760 ;
  LAYER metal1 ;
  RECT 3029.720 178.640 3033.260 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3016.080 178.640 3019.620 179.760 ;
  LAYER metal4 ;
  RECT 3016.080 178.640 3019.620 179.760 ;
  LAYER metal3 ;
  RECT 3016.080 178.640 3019.620 179.760 ;
  LAYER metal2 ;
  RECT 3016.080 178.640 3019.620 179.760 ;
  LAYER metal1 ;
  RECT 3016.080 178.640 3019.620 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3002.440 178.640 3005.980 179.760 ;
  LAYER metal4 ;
  RECT 3002.440 178.640 3005.980 179.760 ;
  LAYER metal3 ;
  RECT 3002.440 178.640 3005.980 179.760 ;
  LAYER metal2 ;
  RECT 3002.440 178.640 3005.980 179.760 ;
  LAYER metal1 ;
  RECT 3002.440 178.640 3005.980 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2989.420 178.640 2992.960 179.760 ;
  LAYER metal4 ;
  RECT 2989.420 178.640 2992.960 179.760 ;
  LAYER metal3 ;
  RECT 2989.420 178.640 2992.960 179.760 ;
  LAYER metal2 ;
  RECT 2989.420 178.640 2992.960 179.760 ;
  LAYER metal1 ;
  RECT 2989.420 178.640 2992.960 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2975.780 178.640 2979.320 179.760 ;
  LAYER metal4 ;
  RECT 2975.780 178.640 2979.320 179.760 ;
  LAYER metal3 ;
  RECT 2975.780 178.640 2979.320 179.760 ;
  LAYER metal2 ;
  RECT 2975.780 178.640 2979.320 179.760 ;
  LAYER metal1 ;
  RECT 2975.780 178.640 2979.320 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2908.200 178.640 2911.740 179.760 ;
  LAYER metal4 ;
  RECT 2908.200 178.640 2911.740 179.760 ;
  LAYER metal3 ;
  RECT 2908.200 178.640 2911.740 179.760 ;
  LAYER metal2 ;
  RECT 2908.200 178.640 2911.740 179.760 ;
  LAYER metal1 ;
  RECT 2908.200 178.640 2911.740 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2895.180 178.640 2898.720 179.760 ;
  LAYER metal4 ;
  RECT 2895.180 178.640 2898.720 179.760 ;
  LAYER metal3 ;
  RECT 2895.180 178.640 2898.720 179.760 ;
  LAYER metal2 ;
  RECT 2895.180 178.640 2898.720 179.760 ;
  LAYER metal1 ;
  RECT 2895.180 178.640 2898.720 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2881.540 178.640 2885.080 179.760 ;
  LAYER metal4 ;
  RECT 2881.540 178.640 2885.080 179.760 ;
  LAYER metal3 ;
  RECT 2881.540 178.640 2885.080 179.760 ;
  LAYER metal2 ;
  RECT 2881.540 178.640 2885.080 179.760 ;
  LAYER metal1 ;
  RECT 2881.540 178.640 2885.080 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2867.900 178.640 2871.440 179.760 ;
  LAYER metal4 ;
  RECT 2867.900 178.640 2871.440 179.760 ;
  LAYER metal3 ;
  RECT 2867.900 178.640 2871.440 179.760 ;
  LAYER metal2 ;
  RECT 2867.900 178.640 2871.440 179.760 ;
  LAYER metal1 ;
  RECT 2867.900 178.640 2871.440 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2854.880 178.640 2858.420 179.760 ;
  LAYER metal4 ;
  RECT 2854.880 178.640 2858.420 179.760 ;
  LAYER metal3 ;
  RECT 2854.880 178.640 2858.420 179.760 ;
  LAYER metal2 ;
  RECT 2854.880 178.640 2858.420 179.760 ;
  LAYER metal1 ;
  RECT 2854.880 178.640 2858.420 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2841.240 178.640 2844.780 179.760 ;
  LAYER metal4 ;
  RECT 2841.240 178.640 2844.780 179.760 ;
  LAYER metal3 ;
  RECT 2841.240 178.640 2844.780 179.760 ;
  LAYER metal2 ;
  RECT 2841.240 178.640 2844.780 179.760 ;
  LAYER metal1 ;
  RECT 2841.240 178.640 2844.780 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2774.280 178.640 2777.820 179.760 ;
  LAYER metal4 ;
  RECT 2774.280 178.640 2777.820 179.760 ;
  LAYER metal3 ;
  RECT 2774.280 178.640 2777.820 179.760 ;
  LAYER metal2 ;
  RECT 2774.280 178.640 2777.820 179.760 ;
  LAYER metal1 ;
  RECT 2774.280 178.640 2777.820 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2760.640 178.640 2764.180 179.760 ;
  LAYER metal4 ;
  RECT 2760.640 178.640 2764.180 179.760 ;
  LAYER metal3 ;
  RECT 2760.640 178.640 2764.180 179.760 ;
  LAYER metal2 ;
  RECT 2760.640 178.640 2764.180 179.760 ;
  LAYER metal1 ;
  RECT 2760.640 178.640 2764.180 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2747.000 178.640 2750.540 179.760 ;
  LAYER metal4 ;
  RECT 2747.000 178.640 2750.540 179.760 ;
  LAYER metal3 ;
  RECT 2747.000 178.640 2750.540 179.760 ;
  LAYER metal2 ;
  RECT 2747.000 178.640 2750.540 179.760 ;
  LAYER metal1 ;
  RECT 2747.000 178.640 2750.540 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2733.980 178.640 2737.520 179.760 ;
  LAYER metal4 ;
  RECT 2733.980 178.640 2737.520 179.760 ;
  LAYER metal3 ;
  RECT 2733.980 178.640 2737.520 179.760 ;
  LAYER metal2 ;
  RECT 2733.980 178.640 2737.520 179.760 ;
  LAYER metal1 ;
  RECT 2733.980 178.640 2737.520 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2720.340 178.640 2723.880 179.760 ;
  LAYER metal4 ;
  RECT 2720.340 178.640 2723.880 179.760 ;
  LAYER metal3 ;
  RECT 2720.340 178.640 2723.880 179.760 ;
  LAYER metal2 ;
  RECT 2720.340 178.640 2723.880 179.760 ;
  LAYER metal1 ;
  RECT 2720.340 178.640 2723.880 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2706.700 178.640 2710.240 179.760 ;
  LAYER metal4 ;
  RECT 2706.700 178.640 2710.240 179.760 ;
  LAYER metal3 ;
  RECT 2706.700 178.640 2710.240 179.760 ;
  LAYER metal2 ;
  RECT 2706.700 178.640 2710.240 179.760 ;
  LAYER metal1 ;
  RECT 2706.700 178.640 2710.240 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2639.740 178.640 2643.280 179.760 ;
  LAYER metal4 ;
  RECT 2639.740 178.640 2643.280 179.760 ;
  LAYER metal3 ;
  RECT 2639.740 178.640 2643.280 179.760 ;
  LAYER metal2 ;
  RECT 2639.740 178.640 2643.280 179.760 ;
  LAYER metal1 ;
  RECT 2639.740 178.640 2643.280 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2626.100 178.640 2629.640 179.760 ;
  LAYER metal4 ;
  RECT 2626.100 178.640 2629.640 179.760 ;
  LAYER metal3 ;
  RECT 2626.100 178.640 2629.640 179.760 ;
  LAYER metal2 ;
  RECT 2626.100 178.640 2629.640 179.760 ;
  LAYER metal1 ;
  RECT 2626.100 178.640 2629.640 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2613.080 178.640 2616.620 179.760 ;
  LAYER metal4 ;
  RECT 2613.080 178.640 2616.620 179.760 ;
  LAYER metal3 ;
  RECT 2613.080 178.640 2616.620 179.760 ;
  LAYER metal2 ;
  RECT 2613.080 178.640 2616.620 179.760 ;
  LAYER metal1 ;
  RECT 2613.080 178.640 2616.620 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2599.440 178.640 2602.980 179.760 ;
  LAYER metal4 ;
  RECT 2599.440 178.640 2602.980 179.760 ;
  LAYER metal3 ;
  RECT 2599.440 178.640 2602.980 179.760 ;
  LAYER metal2 ;
  RECT 2599.440 178.640 2602.980 179.760 ;
  LAYER metal1 ;
  RECT 2599.440 178.640 2602.980 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2585.800 178.640 2589.340 179.760 ;
  LAYER metal4 ;
  RECT 2585.800 178.640 2589.340 179.760 ;
  LAYER metal3 ;
  RECT 2585.800 178.640 2589.340 179.760 ;
  LAYER metal2 ;
  RECT 2585.800 178.640 2589.340 179.760 ;
  LAYER metal1 ;
  RECT 2585.800 178.640 2589.340 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2572.780 178.640 2576.320 179.760 ;
  LAYER metal4 ;
  RECT 2572.780 178.640 2576.320 179.760 ;
  LAYER metal3 ;
  RECT 2572.780 178.640 2576.320 179.760 ;
  LAYER metal2 ;
  RECT 2572.780 178.640 2576.320 179.760 ;
  LAYER metal1 ;
  RECT 2572.780 178.640 2576.320 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2505.200 178.640 2508.740 179.760 ;
  LAYER metal4 ;
  RECT 2505.200 178.640 2508.740 179.760 ;
  LAYER metal3 ;
  RECT 2505.200 178.640 2508.740 179.760 ;
  LAYER metal2 ;
  RECT 2505.200 178.640 2508.740 179.760 ;
  LAYER metal1 ;
  RECT 2505.200 178.640 2508.740 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2491.560 178.640 2495.100 179.760 ;
  LAYER metal4 ;
  RECT 2491.560 178.640 2495.100 179.760 ;
  LAYER metal3 ;
  RECT 2491.560 178.640 2495.100 179.760 ;
  LAYER metal2 ;
  RECT 2491.560 178.640 2495.100 179.760 ;
  LAYER metal1 ;
  RECT 2491.560 178.640 2495.100 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2478.540 178.640 2482.080 179.760 ;
  LAYER metal4 ;
  RECT 2478.540 178.640 2482.080 179.760 ;
  LAYER metal3 ;
  RECT 2478.540 178.640 2482.080 179.760 ;
  LAYER metal2 ;
  RECT 2478.540 178.640 2482.080 179.760 ;
  LAYER metal1 ;
  RECT 2478.540 178.640 2482.080 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2464.900 178.640 2468.440 179.760 ;
  LAYER metal4 ;
  RECT 2464.900 178.640 2468.440 179.760 ;
  LAYER metal3 ;
  RECT 2464.900 178.640 2468.440 179.760 ;
  LAYER metal2 ;
  RECT 2464.900 178.640 2468.440 179.760 ;
  LAYER metal1 ;
  RECT 2464.900 178.640 2468.440 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2451.260 178.640 2454.800 179.760 ;
  LAYER metal4 ;
  RECT 2451.260 178.640 2454.800 179.760 ;
  LAYER metal3 ;
  RECT 2451.260 178.640 2454.800 179.760 ;
  LAYER metal2 ;
  RECT 2451.260 178.640 2454.800 179.760 ;
  LAYER metal1 ;
  RECT 2451.260 178.640 2454.800 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2438.240 178.640 2441.780 179.760 ;
  LAYER metal4 ;
  RECT 2438.240 178.640 2441.780 179.760 ;
  LAYER metal3 ;
  RECT 2438.240 178.640 2441.780 179.760 ;
  LAYER metal2 ;
  RECT 2438.240 178.640 2441.780 179.760 ;
  LAYER metal1 ;
  RECT 2438.240 178.640 2441.780 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2370.660 178.640 2374.200 179.760 ;
  LAYER metal4 ;
  RECT 2370.660 178.640 2374.200 179.760 ;
  LAYER metal3 ;
  RECT 2370.660 178.640 2374.200 179.760 ;
  LAYER metal2 ;
  RECT 2370.660 178.640 2374.200 179.760 ;
  LAYER metal1 ;
  RECT 2370.660 178.640 2374.200 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2357.640 178.640 2361.180 179.760 ;
  LAYER metal4 ;
  RECT 2357.640 178.640 2361.180 179.760 ;
  LAYER metal3 ;
  RECT 2357.640 178.640 2361.180 179.760 ;
  LAYER metal2 ;
  RECT 2357.640 178.640 2361.180 179.760 ;
  LAYER metal1 ;
  RECT 2357.640 178.640 2361.180 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2344.000 178.640 2347.540 179.760 ;
  LAYER metal4 ;
  RECT 2344.000 178.640 2347.540 179.760 ;
  LAYER metal3 ;
  RECT 2344.000 178.640 2347.540 179.760 ;
  LAYER metal2 ;
  RECT 2344.000 178.640 2347.540 179.760 ;
  LAYER metal1 ;
  RECT 2344.000 178.640 2347.540 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2330.360 178.640 2333.900 179.760 ;
  LAYER metal4 ;
  RECT 2330.360 178.640 2333.900 179.760 ;
  LAYER metal3 ;
  RECT 2330.360 178.640 2333.900 179.760 ;
  LAYER metal2 ;
  RECT 2330.360 178.640 2333.900 179.760 ;
  LAYER metal1 ;
  RECT 2330.360 178.640 2333.900 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2317.340 178.640 2320.880 179.760 ;
  LAYER metal4 ;
  RECT 2317.340 178.640 2320.880 179.760 ;
  LAYER metal3 ;
  RECT 2317.340 178.640 2320.880 179.760 ;
  LAYER metal2 ;
  RECT 2317.340 178.640 2320.880 179.760 ;
  LAYER metal1 ;
  RECT 2317.340 178.640 2320.880 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2303.700 178.640 2307.240 179.760 ;
  LAYER metal4 ;
  RECT 2303.700 178.640 2307.240 179.760 ;
  LAYER metal3 ;
  RECT 2303.700 178.640 2307.240 179.760 ;
  LAYER metal2 ;
  RECT 2303.700 178.640 2307.240 179.760 ;
  LAYER metal1 ;
  RECT 2303.700 178.640 2307.240 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2236.740 178.640 2240.280 179.760 ;
  LAYER metal4 ;
  RECT 2236.740 178.640 2240.280 179.760 ;
  LAYER metal3 ;
  RECT 2236.740 178.640 2240.280 179.760 ;
  LAYER metal2 ;
  RECT 2236.740 178.640 2240.280 179.760 ;
  LAYER metal1 ;
  RECT 2236.740 178.640 2240.280 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2223.100 178.640 2226.640 179.760 ;
  LAYER metal4 ;
  RECT 2223.100 178.640 2226.640 179.760 ;
  LAYER metal3 ;
  RECT 2223.100 178.640 2226.640 179.760 ;
  LAYER metal2 ;
  RECT 2223.100 178.640 2226.640 179.760 ;
  LAYER metal1 ;
  RECT 2223.100 178.640 2226.640 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2209.460 178.640 2213.000 179.760 ;
  LAYER metal4 ;
  RECT 2209.460 178.640 2213.000 179.760 ;
  LAYER metal3 ;
  RECT 2209.460 178.640 2213.000 179.760 ;
  LAYER metal2 ;
  RECT 2209.460 178.640 2213.000 179.760 ;
  LAYER metal1 ;
  RECT 2209.460 178.640 2213.000 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2196.440 178.640 2199.980 179.760 ;
  LAYER metal4 ;
  RECT 2196.440 178.640 2199.980 179.760 ;
  LAYER metal3 ;
  RECT 2196.440 178.640 2199.980 179.760 ;
  LAYER metal2 ;
  RECT 2196.440 178.640 2199.980 179.760 ;
  LAYER metal1 ;
  RECT 2196.440 178.640 2199.980 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2182.800 178.640 2186.340 179.760 ;
  LAYER metal4 ;
  RECT 2182.800 178.640 2186.340 179.760 ;
  LAYER metal3 ;
  RECT 2182.800 178.640 2186.340 179.760 ;
  LAYER metal2 ;
  RECT 2182.800 178.640 2186.340 179.760 ;
  LAYER metal1 ;
  RECT 2182.800 178.640 2186.340 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2169.160 178.640 2172.700 179.760 ;
  LAYER metal4 ;
  RECT 2169.160 178.640 2172.700 179.760 ;
  LAYER metal3 ;
  RECT 2169.160 178.640 2172.700 179.760 ;
  LAYER metal2 ;
  RECT 2169.160 178.640 2172.700 179.760 ;
  LAYER metal1 ;
  RECT 2169.160 178.640 2172.700 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2102.200 178.640 2105.740 179.760 ;
  LAYER metal4 ;
  RECT 2102.200 178.640 2105.740 179.760 ;
  LAYER metal3 ;
  RECT 2102.200 178.640 2105.740 179.760 ;
  LAYER metal2 ;
  RECT 2102.200 178.640 2105.740 179.760 ;
  LAYER metal1 ;
  RECT 2102.200 178.640 2105.740 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2088.560 178.640 2092.100 179.760 ;
  LAYER metal4 ;
  RECT 2088.560 178.640 2092.100 179.760 ;
  LAYER metal3 ;
  RECT 2088.560 178.640 2092.100 179.760 ;
  LAYER metal2 ;
  RECT 2088.560 178.640 2092.100 179.760 ;
  LAYER metal1 ;
  RECT 2088.560 178.640 2092.100 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2074.920 178.640 2078.460 179.760 ;
  LAYER metal4 ;
  RECT 2074.920 178.640 2078.460 179.760 ;
  LAYER metal3 ;
  RECT 2074.920 178.640 2078.460 179.760 ;
  LAYER metal2 ;
  RECT 2074.920 178.640 2078.460 179.760 ;
  LAYER metal1 ;
  RECT 2074.920 178.640 2078.460 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2061.900 178.640 2065.440 179.760 ;
  LAYER metal4 ;
  RECT 2061.900 178.640 2065.440 179.760 ;
  LAYER metal3 ;
  RECT 2061.900 178.640 2065.440 179.760 ;
  LAYER metal2 ;
  RECT 2061.900 178.640 2065.440 179.760 ;
  LAYER metal1 ;
  RECT 2061.900 178.640 2065.440 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2048.260 178.640 2051.800 179.760 ;
  LAYER metal4 ;
  RECT 2048.260 178.640 2051.800 179.760 ;
  LAYER metal3 ;
  RECT 2048.260 178.640 2051.800 179.760 ;
  LAYER metal2 ;
  RECT 2048.260 178.640 2051.800 179.760 ;
  LAYER metal1 ;
  RECT 2048.260 178.640 2051.800 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2034.620 178.640 2038.160 179.760 ;
  LAYER metal4 ;
  RECT 2034.620 178.640 2038.160 179.760 ;
  LAYER metal3 ;
  RECT 2034.620 178.640 2038.160 179.760 ;
  LAYER metal2 ;
  RECT 2034.620 178.640 2038.160 179.760 ;
  LAYER metal1 ;
  RECT 2034.620 178.640 2038.160 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1967.660 178.640 1971.200 179.760 ;
  LAYER metal4 ;
  RECT 1967.660 178.640 1971.200 179.760 ;
  LAYER metal3 ;
  RECT 1967.660 178.640 1971.200 179.760 ;
  LAYER metal2 ;
  RECT 1967.660 178.640 1971.200 179.760 ;
  LAYER metal1 ;
  RECT 1967.660 178.640 1971.200 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1954.020 178.640 1957.560 179.760 ;
  LAYER metal4 ;
  RECT 1954.020 178.640 1957.560 179.760 ;
  LAYER metal3 ;
  RECT 1954.020 178.640 1957.560 179.760 ;
  LAYER metal2 ;
  RECT 1954.020 178.640 1957.560 179.760 ;
  LAYER metal1 ;
  RECT 1954.020 178.640 1957.560 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1941.000 178.640 1944.540 179.760 ;
  LAYER metal4 ;
  RECT 1941.000 178.640 1944.540 179.760 ;
  LAYER metal3 ;
  RECT 1941.000 178.640 1944.540 179.760 ;
  LAYER metal2 ;
  RECT 1941.000 178.640 1944.540 179.760 ;
  LAYER metal1 ;
  RECT 1941.000 178.640 1944.540 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1927.360 178.640 1930.900 179.760 ;
  LAYER metal4 ;
  RECT 1927.360 178.640 1930.900 179.760 ;
  LAYER metal3 ;
  RECT 1927.360 178.640 1930.900 179.760 ;
  LAYER metal2 ;
  RECT 1927.360 178.640 1930.900 179.760 ;
  LAYER metal1 ;
  RECT 1927.360 178.640 1930.900 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1913.720 178.640 1917.260 179.760 ;
  LAYER metal4 ;
  RECT 1913.720 178.640 1917.260 179.760 ;
  LAYER metal3 ;
  RECT 1913.720 178.640 1917.260 179.760 ;
  LAYER metal2 ;
  RECT 1913.720 178.640 1917.260 179.760 ;
  LAYER metal1 ;
  RECT 1913.720 178.640 1917.260 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1900.700 178.640 1904.240 179.760 ;
  LAYER metal4 ;
  RECT 1900.700 178.640 1904.240 179.760 ;
  LAYER metal3 ;
  RECT 1900.700 178.640 1904.240 179.760 ;
  LAYER metal2 ;
  RECT 1900.700 178.640 1904.240 179.760 ;
  LAYER metal1 ;
  RECT 1900.700 178.640 1904.240 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1833.120 178.640 1836.660 179.760 ;
  LAYER metal4 ;
  RECT 1833.120 178.640 1836.660 179.760 ;
  LAYER metal3 ;
  RECT 1833.120 178.640 1836.660 179.760 ;
  LAYER metal2 ;
  RECT 1833.120 178.640 1836.660 179.760 ;
  LAYER metal1 ;
  RECT 1833.120 178.640 1836.660 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1821.960 178.640 1825.500 179.760 ;
  LAYER metal4 ;
  RECT 1821.960 178.640 1825.500 179.760 ;
  LAYER metal3 ;
  RECT 1821.960 178.640 1825.500 179.760 ;
  LAYER metal2 ;
  RECT 1821.960 178.640 1825.500 179.760 ;
  LAYER metal1 ;
  RECT 1821.960 178.640 1825.500 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1805.840 178.640 1809.380 179.760 ;
  LAYER metal4 ;
  RECT 1805.840 178.640 1809.380 179.760 ;
  LAYER metal3 ;
  RECT 1805.840 178.640 1809.380 179.760 ;
  LAYER metal2 ;
  RECT 1805.840 178.640 1809.380 179.760 ;
  LAYER metal1 ;
  RECT 1805.840 178.640 1809.380 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1797.160 178.640 1800.700 179.760 ;
  LAYER metal4 ;
  RECT 1797.160 178.640 1800.700 179.760 ;
  LAYER metal3 ;
  RECT 1797.160 178.640 1800.700 179.760 ;
  LAYER metal2 ;
  RECT 1797.160 178.640 1800.700 179.760 ;
  LAYER metal1 ;
  RECT 1797.160 178.640 1800.700 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1784.140 178.640 1787.680 179.760 ;
  LAYER metal4 ;
  RECT 1784.140 178.640 1787.680 179.760 ;
  LAYER metal3 ;
  RECT 1784.140 178.640 1787.680 179.760 ;
  LAYER metal2 ;
  RECT 1784.140 178.640 1787.680 179.760 ;
  LAYER metal1 ;
  RECT 1784.140 178.640 1787.680 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1771.120 178.640 1774.660 179.760 ;
  LAYER metal4 ;
  RECT 1771.120 178.640 1774.660 179.760 ;
  LAYER metal3 ;
  RECT 1771.120 178.640 1774.660 179.760 ;
  LAYER metal2 ;
  RECT 1771.120 178.640 1774.660 179.760 ;
  LAYER metal1 ;
  RECT 1771.120 178.640 1774.660 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1685.560 178.640 1689.100 179.760 ;
  LAYER metal4 ;
  RECT 1685.560 178.640 1689.100 179.760 ;
  LAYER metal3 ;
  RECT 1685.560 178.640 1689.100 179.760 ;
  LAYER metal2 ;
  RECT 1685.560 178.640 1689.100 179.760 ;
  LAYER metal1 ;
  RECT 1685.560 178.640 1689.100 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1672.540 178.640 1676.080 179.760 ;
  LAYER metal4 ;
  RECT 1672.540 178.640 1676.080 179.760 ;
  LAYER metal3 ;
  RECT 1672.540 178.640 1676.080 179.760 ;
  LAYER metal2 ;
  RECT 1672.540 178.640 1676.080 179.760 ;
  LAYER metal1 ;
  RECT 1672.540 178.640 1676.080 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1658.900 178.640 1662.440 179.760 ;
  LAYER metal4 ;
  RECT 1658.900 178.640 1662.440 179.760 ;
  LAYER metal3 ;
  RECT 1658.900 178.640 1662.440 179.760 ;
  LAYER metal2 ;
  RECT 1658.900 178.640 1662.440 179.760 ;
  LAYER metal1 ;
  RECT 1658.900 178.640 1662.440 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1645.260 178.640 1648.800 179.760 ;
  LAYER metal4 ;
  RECT 1645.260 178.640 1648.800 179.760 ;
  LAYER metal3 ;
  RECT 1645.260 178.640 1648.800 179.760 ;
  LAYER metal2 ;
  RECT 1645.260 178.640 1648.800 179.760 ;
  LAYER metal1 ;
  RECT 1645.260 178.640 1648.800 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1632.240 178.640 1635.780 179.760 ;
  LAYER metal4 ;
  RECT 1632.240 178.640 1635.780 179.760 ;
  LAYER metal3 ;
  RECT 1632.240 178.640 1635.780 179.760 ;
  LAYER metal2 ;
  RECT 1632.240 178.640 1635.780 179.760 ;
  LAYER metal1 ;
  RECT 1632.240 178.640 1635.780 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1618.600 178.640 1622.140 179.760 ;
  LAYER metal4 ;
  RECT 1618.600 178.640 1622.140 179.760 ;
  LAYER metal3 ;
  RECT 1618.600 178.640 1622.140 179.760 ;
  LAYER metal2 ;
  RECT 1618.600 178.640 1622.140 179.760 ;
  LAYER metal1 ;
  RECT 1618.600 178.640 1622.140 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1551.640 178.640 1555.180 179.760 ;
  LAYER metal4 ;
  RECT 1551.640 178.640 1555.180 179.760 ;
  LAYER metal3 ;
  RECT 1551.640 178.640 1555.180 179.760 ;
  LAYER metal2 ;
  RECT 1551.640 178.640 1555.180 179.760 ;
  LAYER metal1 ;
  RECT 1551.640 178.640 1555.180 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1538.000 178.640 1541.540 179.760 ;
  LAYER metal4 ;
  RECT 1538.000 178.640 1541.540 179.760 ;
  LAYER metal3 ;
  RECT 1538.000 178.640 1541.540 179.760 ;
  LAYER metal2 ;
  RECT 1538.000 178.640 1541.540 179.760 ;
  LAYER metal1 ;
  RECT 1538.000 178.640 1541.540 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1524.360 178.640 1527.900 179.760 ;
  LAYER metal4 ;
  RECT 1524.360 178.640 1527.900 179.760 ;
  LAYER metal3 ;
  RECT 1524.360 178.640 1527.900 179.760 ;
  LAYER metal2 ;
  RECT 1524.360 178.640 1527.900 179.760 ;
  LAYER metal1 ;
  RECT 1524.360 178.640 1527.900 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1511.340 178.640 1514.880 179.760 ;
  LAYER metal4 ;
  RECT 1511.340 178.640 1514.880 179.760 ;
  LAYER metal3 ;
  RECT 1511.340 178.640 1514.880 179.760 ;
  LAYER metal2 ;
  RECT 1511.340 178.640 1514.880 179.760 ;
  LAYER metal1 ;
  RECT 1511.340 178.640 1514.880 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1497.700 178.640 1501.240 179.760 ;
  LAYER metal4 ;
  RECT 1497.700 178.640 1501.240 179.760 ;
  LAYER metal3 ;
  RECT 1497.700 178.640 1501.240 179.760 ;
  LAYER metal2 ;
  RECT 1497.700 178.640 1501.240 179.760 ;
  LAYER metal1 ;
  RECT 1497.700 178.640 1501.240 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1484.060 178.640 1487.600 179.760 ;
  LAYER metal4 ;
  RECT 1484.060 178.640 1487.600 179.760 ;
  LAYER metal3 ;
  RECT 1484.060 178.640 1487.600 179.760 ;
  LAYER metal2 ;
  RECT 1484.060 178.640 1487.600 179.760 ;
  LAYER metal1 ;
  RECT 1484.060 178.640 1487.600 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1417.100 178.640 1420.640 179.760 ;
  LAYER metal4 ;
  RECT 1417.100 178.640 1420.640 179.760 ;
  LAYER metal3 ;
  RECT 1417.100 178.640 1420.640 179.760 ;
  LAYER metal2 ;
  RECT 1417.100 178.640 1420.640 179.760 ;
  LAYER metal1 ;
  RECT 1417.100 178.640 1420.640 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1403.460 178.640 1407.000 179.760 ;
  LAYER metal4 ;
  RECT 1403.460 178.640 1407.000 179.760 ;
  LAYER metal3 ;
  RECT 1403.460 178.640 1407.000 179.760 ;
  LAYER metal2 ;
  RECT 1403.460 178.640 1407.000 179.760 ;
  LAYER metal1 ;
  RECT 1403.460 178.640 1407.000 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1390.440 178.640 1393.980 179.760 ;
  LAYER metal4 ;
  RECT 1390.440 178.640 1393.980 179.760 ;
  LAYER metal3 ;
  RECT 1390.440 178.640 1393.980 179.760 ;
  LAYER metal2 ;
  RECT 1390.440 178.640 1393.980 179.760 ;
  LAYER metal1 ;
  RECT 1390.440 178.640 1393.980 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1376.800 178.640 1380.340 179.760 ;
  LAYER metal4 ;
  RECT 1376.800 178.640 1380.340 179.760 ;
  LAYER metal3 ;
  RECT 1376.800 178.640 1380.340 179.760 ;
  LAYER metal2 ;
  RECT 1376.800 178.640 1380.340 179.760 ;
  LAYER metal1 ;
  RECT 1376.800 178.640 1380.340 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1363.160 178.640 1366.700 179.760 ;
  LAYER metal4 ;
  RECT 1363.160 178.640 1366.700 179.760 ;
  LAYER metal3 ;
  RECT 1363.160 178.640 1366.700 179.760 ;
  LAYER metal2 ;
  RECT 1363.160 178.640 1366.700 179.760 ;
  LAYER metal1 ;
  RECT 1363.160 178.640 1366.700 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1350.140 178.640 1353.680 179.760 ;
  LAYER metal4 ;
  RECT 1350.140 178.640 1353.680 179.760 ;
  LAYER metal3 ;
  RECT 1350.140 178.640 1353.680 179.760 ;
  LAYER metal2 ;
  RECT 1350.140 178.640 1353.680 179.760 ;
  LAYER metal1 ;
  RECT 1350.140 178.640 1353.680 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1282.560 178.640 1286.100 179.760 ;
  LAYER metal4 ;
  RECT 1282.560 178.640 1286.100 179.760 ;
  LAYER metal3 ;
  RECT 1282.560 178.640 1286.100 179.760 ;
  LAYER metal2 ;
  RECT 1282.560 178.640 1286.100 179.760 ;
  LAYER metal1 ;
  RECT 1282.560 178.640 1286.100 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1268.920 178.640 1272.460 179.760 ;
  LAYER metal4 ;
  RECT 1268.920 178.640 1272.460 179.760 ;
  LAYER metal3 ;
  RECT 1268.920 178.640 1272.460 179.760 ;
  LAYER metal2 ;
  RECT 1268.920 178.640 1272.460 179.760 ;
  LAYER metal1 ;
  RECT 1268.920 178.640 1272.460 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1255.900 178.640 1259.440 179.760 ;
  LAYER metal4 ;
  RECT 1255.900 178.640 1259.440 179.760 ;
  LAYER metal3 ;
  RECT 1255.900 178.640 1259.440 179.760 ;
  LAYER metal2 ;
  RECT 1255.900 178.640 1259.440 179.760 ;
  LAYER metal1 ;
  RECT 1255.900 178.640 1259.440 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1242.260 178.640 1245.800 179.760 ;
  LAYER metal4 ;
  RECT 1242.260 178.640 1245.800 179.760 ;
  LAYER metal3 ;
  RECT 1242.260 178.640 1245.800 179.760 ;
  LAYER metal2 ;
  RECT 1242.260 178.640 1245.800 179.760 ;
  LAYER metal1 ;
  RECT 1242.260 178.640 1245.800 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1228.620 178.640 1232.160 179.760 ;
  LAYER metal4 ;
  RECT 1228.620 178.640 1232.160 179.760 ;
  LAYER metal3 ;
  RECT 1228.620 178.640 1232.160 179.760 ;
  LAYER metal2 ;
  RECT 1228.620 178.640 1232.160 179.760 ;
  LAYER metal1 ;
  RECT 1228.620 178.640 1232.160 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1215.600 178.640 1219.140 179.760 ;
  LAYER metal4 ;
  RECT 1215.600 178.640 1219.140 179.760 ;
  LAYER metal3 ;
  RECT 1215.600 178.640 1219.140 179.760 ;
  LAYER metal2 ;
  RECT 1215.600 178.640 1219.140 179.760 ;
  LAYER metal1 ;
  RECT 1215.600 178.640 1219.140 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1148.020 178.640 1151.560 179.760 ;
  LAYER metal4 ;
  RECT 1148.020 178.640 1151.560 179.760 ;
  LAYER metal3 ;
  RECT 1148.020 178.640 1151.560 179.760 ;
  LAYER metal2 ;
  RECT 1148.020 178.640 1151.560 179.760 ;
  LAYER metal1 ;
  RECT 1148.020 178.640 1151.560 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1135.000 178.640 1138.540 179.760 ;
  LAYER metal4 ;
  RECT 1135.000 178.640 1138.540 179.760 ;
  LAYER metal3 ;
  RECT 1135.000 178.640 1138.540 179.760 ;
  LAYER metal2 ;
  RECT 1135.000 178.640 1138.540 179.760 ;
  LAYER metal1 ;
  RECT 1135.000 178.640 1138.540 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1121.360 178.640 1124.900 179.760 ;
  LAYER metal4 ;
  RECT 1121.360 178.640 1124.900 179.760 ;
  LAYER metal3 ;
  RECT 1121.360 178.640 1124.900 179.760 ;
  LAYER metal2 ;
  RECT 1121.360 178.640 1124.900 179.760 ;
  LAYER metal1 ;
  RECT 1121.360 178.640 1124.900 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1107.720 178.640 1111.260 179.760 ;
  LAYER metal4 ;
  RECT 1107.720 178.640 1111.260 179.760 ;
  LAYER metal3 ;
  RECT 1107.720 178.640 1111.260 179.760 ;
  LAYER metal2 ;
  RECT 1107.720 178.640 1111.260 179.760 ;
  LAYER metal1 ;
  RECT 1107.720 178.640 1111.260 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1094.700 178.640 1098.240 179.760 ;
  LAYER metal4 ;
  RECT 1094.700 178.640 1098.240 179.760 ;
  LAYER metal3 ;
  RECT 1094.700 178.640 1098.240 179.760 ;
  LAYER metal2 ;
  RECT 1094.700 178.640 1098.240 179.760 ;
  LAYER metal1 ;
  RECT 1094.700 178.640 1098.240 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1081.060 178.640 1084.600 179.760 ;
  LAYER metal4 ;
  RECT 1081.060 178.640 1084.600 179.760 ;
  LAYER metal3 ;
  RECT 1081.060 178.640 1084.600 179.760 ;
  LAYER metal2 ;
  RECT 1081.060 178.640 1084.600 179.760 ;
  LAYER metal1 ;
  RECT 1081.060 178.640 1084.600 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1014.100 178.640 1017.640 179.760 ;
  LAYER metal4 ;
  RECT 1014.100 178.640 1017.640 179.760 ;
  LAYER metal3 ;
  RECT 1014.100 178.640 1017.640 179.760 ;
  LAYER metal2 ;
  RECT 1014.100 178.640 1017.640 179.760 ;
  LAYER metal1 ;
  RECT 1014.100 178.640 1017.640 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1000.460 178.640 1004.000 179.760 ;
  LAYER metal4 ;
  RECT 1000.460 178.640 1004.000 179.760 ;
  LAYER metal3 ;
  RECT 1000.460 178.640 1004.000 179.760 ;
  LAYER metal2 ;
  RECT 1000.460 178.640 1004.000 179.760 ;
  LAYER metal1 ;
  RECT 1000.460 178.640 1004.000 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 986.820 178.640 990.360 179.760 ;
  LAYER metal4 ;
  RECT 986.820 178.640 990.360 179.760 ;
  LAYER metal3 ;
  RECT 986.820 178.640 990.360 179.760 ;
  LAYER metal2 ;
  RECT 986.820 178.640 990.360 179.760 ;
  LAYER metal1 ;
  RECT 986.820 178.640 990.360 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 973.800 178.640 977.340 179.760 ;
  LAYER metal4 ;
  RECT 973.800 178.640 977.340 179.760 ;
  LAYER metal3 ;
  RECT 973.800 178.640 977.340 179.760 ;
  LAYER metal2 ;
  RECT 973.800 178.640 977.340 179.760 ;
  LAYER metal1 ;
  RECT 973.800 178.640 977.340 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 960.160 178.640 963.700 179.760 ;
  LAYER metal4 ;
  RECT 960.160 178.640 963.700 179.760 ;
  LAYER metal3 ;
  RECT 960.160 178.640 963.700 179.760 ;
  LAYER metal2 ;
  RECT 960.160 178.640 963.700 179.760 ;
  LAYER metal1 ;
  RECT 960.160 178.640 963.700 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 946.520 178.640 950.060 179.760 ;
  LAYER metal4 ;
  RECT 946.520 178.640 950.060 179.760 ;
  LAYER metal3 ;
  RECT 946.520 178.640 950.060 179.760 ;
  LAYER metal2 ;
  RECT 946.520 178.640 950.060 179.760 ;
  LAYER metal1 ;
  RECT 946.520 178.640 950.060 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 881.420 178.640 884.960 179.760 ;
  LAYER metal4 ;
  RECT 881.420 178.640 884.960 179.760 ;
  LAYER metal3 ;
  RECT 881.420 178.640 884.960 179.760 ;
  LAYER metal2 ;
  RECT 881.420 178.640 884.960 179.760 ;
  LAYER metal1 ;
  RECT 881.420 178.640 884.960 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 865.920 178.640 869.460 179.760 ;
  LAYER metal4 ;
  RECT 865.920 178.640 869.460 179.760 ;
  LAYER metal3 ;
  RECT 865.920 178.640 869.460 179.760 ;
  LAYER metal2 ;
  RECT 865.920 178.640 869.460 179.760 ;
  LAYER metal1 ;
  RECT 865.920 178.640 869.460 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 852.280 178.640 855.820 179.760 ;
  LAYER metal4 ;
  RECT 852.280 178.640 855.820 179.760 ;
  LAYER metal3 ;
  RECT 852.280 178.640 855.820 179.760 ;
  LAYER metal2 ;
  RECT 852.280 178.640 855.820 179.760 ;
  LAYER metal1 ;
  RECT 852.280 178.640 855.820 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 839.260 178.640 842.800 179.760 ;
  LAYER metal4 ;
  RECT 839.260 178.640 842.800 179.760 ;
  LAYER metal3 ;
  RECT 839.260 178.640 842.800 179.760 ;
  LAYER metal2 ;
  RECT 839.260 178.640 842.800 179.760 ;
  LAYER metal1 ;
  RECT 839.260 178.640 842.800 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 825.620 178.640 829.160 179.760 ;
  LAYER metal4 ;
  RECT 825.620 178.640 829.160 179.760 ;
  LAYER metal3 ;
  RECT 825.620 178.640 829.160 179.760 ;
  LAYER metal2 ;
  RECT 825.620 178.640 829.160 179.760 ;
  LAYER metal1 ;
  RECT 825.620 178.640 829.160 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 811.980 178.640 815.520 179.760 ;
  LAYER metal4 ;
  RECT 811.980 178.640 815.520 179.760 ;
  LAYER metal3 ;
  RECT 811.980 178.640 815.520 179.760 ;
  LAYER metal2 ;
  RECT 811.980 178.640 815.520 179.760 ;
  LAYER metal1 ;
  RECT 811.980 178.640 815.520 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 745.020 178.640 748.560 179.760 ;
  LAYER metal4 ;
  RECT 745.020 178.640 748.560 179.760 ;
  LAYER metal3 ;
  RECT 745.020 178.640 748.560 179.760 ;
  LAYER metal2 ;
  RECT 745.020 178.640 748.560 179.760 ;
  LAYER metal1 ;
  RECT 745.020 178.640 748.560 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 731.380 178.640 734.920 179.760 ;
  LAYER metal4 ;
  RECT 731.380 178.640 734.920 179.760 ;
  LAYER metal3 ;
  RECT 731.380 178.640 734.920 179.760 ;
  LAYER metal2 ;
  RECT 731.380 178.640 734.920 179.760 ;
  LAYER metal1 ;
  RECT 731.380 178.640 734.920 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 718.360 178.640 721.900 179.760 ;
  LAYER metal4 ;
  RECT 718.360 178.640 721.900 179.760 ;
  LAYER metal3 ;
  RECT 718.360 178.640 721.900 179.760 ;
  LAYER metal2 ;
  RECT 718.360 178.640 721.900 179.760 ;
  LAYER metal1 ;
  RECT 718.360 178.640 721.900 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 704.720 178.640 708.260 179.760 ;
  LAYER metal4 ;
  RECT 704.720 178.640 708.260 179.760 ;
  LAYER metal3 ;
  RECT 704.720 178.640 708.260 179.760 ;
  LAYER metal2 ;
  RECT 704.720 178.640 708.260 179.760 ;
  LAYER metal1 ;
  RECT 704.720 178.640 708.260 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 691.080 178.640 694.620 179.760 ;
  LAYER metal4 ;
  RECT 691.080 178.640 694.620 179.760 ;
  LAYER metal3 ;
  RECT 691.080 178.640 694.620 179.760 ;
  LAYER metal2 ;
  RECT 691.080 178.640 694.620 179.760 ;
  LAYER metal1 ;
  RECT 691.080 178.640 694.620 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 678.060 178.640 681.600 179.760 ;
  LAYER metal4 ;
  RECT 678.060 178.640 681.600 179.760 ;
  LAYER metal3 ;
  RECT 678.060 178.640 681.600 179.760 ;
  LAYER metal2 ;
  RECT 678.060 178.640 681.600 179.760 ;
  LAYER metal1 ;
  RECT 678.060 178.640 681.600 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 610.480 178.640 614.020 179.760 ;
  LAYER metal4 ;
  RECT 610.480 178.640 614.020 179.760 ;
  LAYER metal3 ;
  RECT 610.480 178.640 614.020 179.760 ;
  LAYER metal2 ;
  RECT 610.480 178.640 614.020 179.760 ;
  LAYER metal1 ;
  RECT 610.480 178.640 614.020 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 597.460 178.640 601.000 179.760 ;
  LAYER metal4 ;
  RECT 597.460 178.640 601.000 179.760 ;
  LAYER metal3 ;
  RECT 597.460 178.640 601.000 179.760 ;
  LAYER metal2 ;
  RECT 597.460 178.640 601.000 179.760 ;
  LAYER metal1 ;
  RECT 597.460 178.640 601.000 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 583.820 178.640 587.360 179.760 ;
  LAYER metal4 ;
  RECT 583.820 178.640 587.360 179.760 ;
  LAYER metal3 ;
  RECT 583.820 178.640 587.360 179.760 ;
  LAYER metal2 ;
  RECT 583.820 178.640 587.360 179.760 ;
  LAYER metal1 ;
  RECT 583.820 178.640 587.360 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 570.180 178.640 573.720 179.760 ;
  LAYER metal4 ;
  RECT 570.180 178.640 573.720 179.760 ;
  LAYER metal3 ;
  RECT 570.180 178.640 573.720 179.760 ;
  LAYER metal2 ;
  RECT 570.180 178.640 573.720 179.760 ;
  LAYER metal1 ;
  RECT 570.180 178.640 573.720 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 557.160 178.640 560.700 179.760 ;
  LAYER metal4 ;
  RECT 557.160 178.640 560.700 179.760 ;
  LAYER metal3 ;
  RECT 557.160 178.640 560.700 179.760 ;
  LAYER metal2 ;
  RECT 557.160 178.640 560.700 179.760 ;
  LAYER metal1 ;
  RECT 557.160 178.640 560.700 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 543.520 178.640 547.060 179.760 ;
  LAYER metal4 ;
  RECT 543.520 178.640 547.060 179.760 ;
  LAYER metal3 ;
  RECT 543.520 178.640 547.060 179.760 ;
  LAYER metal2 ;
  RECT 543.520 178.640 547.060 179.760 ;
  LAYER metal1 ;
  RECT 543.520 178.640 547.060 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 475.940 178.640 479.480 179.760 ;
  LAYER metal4 ;
  RECT 475.940 178.640 479.480 179.760 ;
  LAYER metal3 ;
  RECT 475.940 178.640 479.480 179.760 ;
  LAYER metal2 ;
  RECT 475.940 178.640 479.480 179.760 ;
  LAYER metal1 ;
  RECT 475.940 178.640 479.480 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 462.920 178.640 466.460 179.760 ;
  LAYER metal4 ;
  RECT 462.920 178.640 466.460 179.760 ;
  LAYER metal3 ;
  RECT 462.920 178.640 466.460 179.760 ;
  LAYER metal2 ;
  RECT 462.920 178.640 466.460 179.760 ;
  LAYER metal1 ;
  RECT 462.920 178.640 466.460 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 451.760 178.640 455.300 179.760 ;
  LAYER metal4 ;
  RECT 451.760 178.640 455.300 179.760 ;
  LAYER metal3 ;
  RECT 451.760 178.640 455.300 179.760 ;
  LAYER metal2 ;
  RECT 451.760 178.640 455.300 179.760 ;
  LAYER metal1 ;
  RECT 451.760 178.640 455.300 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 435.640 178.640 439.180 179.760 ;
  LAYER metal4 ;
  RECT 435.640 178.640 439.180 179.760 ;
  LAYER metal3 ;
  RECT 435.640 178.640 439.180 179.760 ;
  LAYER metal2 ;
  RECT 435.640 178.640 439.180 179.760 ;
  LAYER metal1 ;
  RECT 435.640 178.640 439.180 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 422.620 178.640 426.160 179.760 ;
  LAYER metal4 ;
  RECT 422.620 178.640 426.160 179.760 ;
  LAYER metal3 ;
  RECT 422.620 178.640 426.160 179.760 ;
  LAYER metal2 ;
  RECT 422.620 178.640 426.160 179.760 ;
  LAYER metal1 ;
  RECT 422.620 178.640 426.160 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 408.980 178.640 412.520 179.760 ;
  LAYER metal4 ;
  RECT 408.980 178.640 412.520 179.760 ;
  LAYER metal3 ;
  RECT 408.980 178.640 412.520 179.760 ;
  LAYER metal2 ;
  RECT 408.980 178.640 412.520 179.760 ;
  LAYER metal1 ;
  RECT 408.980 178.640 412.520 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 342.020 178.640 345.560 179.760 ;
  LAYER metal4 ;
  RECT 342.020 178.640 345.560 179.760 ;
  LAYER metal3 ;
  RECT 342.020 178.640 345.560 179.760 ;
  LAYER metal2 ;
  RECT 342.020 178.640 345.560 179.760 ;
  LAYER metal1 ;
  RECT 342.020 178.640 345.560 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 328.380 178.640 331.920 179.760 ;
  LAYER metal4 ;
  RECT 328.380 178.640 331.920 179.760 ;
  LAYER metal3 ;
  RECT 328.380 178.640 331.920 179.760 ;
  LAYER metal2 ;
  RECT 328.380 178.640 331.920 179.760 ;
  LAYER metal1 ;
  RECT 328.380 178.640 331.920 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 314.740 178.640 318.280 179.760 ;
  LAYER metal4 ;
  RECT 314.740 178.640 318.280 179.760 ;
  LAYER metal3 ;
  RECT 314.740 178.640 318.280 179.760 ;
  LAYER metal2 ;
  RECT 314.740 178.640 318.280 179.760 ;
  LAYER metal1 ;
  RECT 314.740 178.640 318.280 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 301.720 178.640 305.260 179.760 ;
  LAYER metal4 ;
  RECT 301.720 178.640 305.260 179.760 ;
  LAYER metal3 ;
  RECT 301.720 178.640 305.260 179.760 ;
  LAYER metal2 ;
  RECT 301.720 178.640 305.260 179.760 ;
  LAYER metal1 ;
  RECT 301.720 178.640 305.260 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 288.080 178.640 291.620 179.760 ;
  LAYER metal4 ;
  RECT 288.080 178.640 291.620 179.760 ;
  LAYER metal3 ;
  RECT 288.080 178.640 291.620 179.760 ;
  LAYER metal2 ;
  RECT 288.080 178.640 291.620 179.760 ;
  LAYER metal1 ;
  RECT 288.080 178.640 291.620 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 274.440 178.640 277.980 179.760 ;
  LAYER metal4 ;
  RECT 274.440 178.640 277.980 179.760 ;
  LAYER metal3 ;
  RECT 274.440 178.640 277.980 179.760 ;
  LAYER metal2 ;
  RECT 274.440 178.640 277.980 179.760 ;
  LAYER metal1 ;
  RECT 274.440 178.640 277.980 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 207.480 178.640 211.020 179.760 ;
  LAYER metal4 ;
  RECT 207.480 178.640 211.020 179.760 ;
  LAYER metal3 ;
  RECT 207.480 178.640 211.020 179.760 ;
  LAYER metal2 ;
  RECT 207.480 178.640 211.020 179.760 ;
  LAYER metal1 ;
  RECT 207.480 178.640 211.020 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 193.840 178.640 197.380 179.760 ;
  LAYER metal4 ;
  RECT 193.840 178.640 197.380 179.760 ;
  LAYER metal3 ;
  RECT 193.840 178.640 197.380 179.760 ;
  LAYER metal2 ;
  RECT 193.840 178.640 197.380 179.760 ;
  LAYER metal1 ;
  RECT 193.840 178.640 197.380 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 180.820 178.640 184.360 179.760 ;
  LAYER metal4 ;
  RECT 180.820 178.640 184.360 179.760 ;
  LAYER metal3 ;
  RECT 180.820 178.640 184.360 179.760 ;
  LAYER metal2 ;
  RECT 180.820 178.640 184.360 179.760 ;
  LAYER metal1 ;
  RECT 180.820 178.640 184.360 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 167.180 178.640 170.720 179.760 ;
  LAYER metal4 ;
  RECT 167.180 178.640 170.720 179.760 ;
  LAYER metal3 ;
  RECT 167.180 178.640 170.720 179.760 ;
  LAYER metal2 ;
  RECT 167.180 178.640 170.720 179.760 ;
  LAYER metal1 ;
  RECT 167.180 178.640 170.720 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 153.540 178.640 157.080 179.760 ;
  LAYER metal4 ;
  RECT 153.540 178.640 157.080 179.760 ;
  LAYER metal3 ;
  RECT 153.540 178.640 157.080 179.760 ;
  LAYER metal2 ;
  RECT 153.540 178.640 157.080 179.760 ;
  LAYER metal1 ;
  RECT 153.540 178.640 157.080 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 140.520 178.640 144.060 179.760 ;
  LAYER metal4 ;
  RECT 140.520 178.640 144.060 179.760 ;
  LAYER metal3 ;
  RECT 140.520 178.640 144.060 179.760 ;
  LAYER metal2 ;
  RECT 140.520 178.640 144.060 179.760 ;
  LAYER metal1 ;
  RECT 140.520 178.640 144.060 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 72.940 178.640 76.480 179.760 ;
  LAYER metal4 ;
  RECT 72.940 178.640 76.480 179.760 ;
  LAYER metal3 ;
  RECT 72.940 178.640 76.480 179.760 ;
  LAYER metal2 ;
  RECT 72.940 178.640 76.480 179.760 ;
  LAYER metal1 ;
  RECT 72.940 178.640 76.480 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 59.300 178.640 62.840 179.760 ;
  LAYER metal4 ;
  RECT 59.300 178.640 62.840 179.760 ;
  LAYER metal3 ;
  RECT 59.300 178.640 62.840 179.760 ;
  LAYER metal2 ;
  RECT 59.300 178.640 62.840 179.760 ;
  LAYER metal1 ;
  RECT 59.300 178.640 62.840 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 46.280 178.640 49.820 179.760 ;
  LAYER metal4 ;
  RECT 46.280 178.640 49.820 179.760 ;
  LAYER metal3 ;
  RECT 46.280 178.640 49.820 179.760 ;
  LAYER metal2 ;
  RECT 46.280 178.640 49.820 179.760 ;
  LAYER metal1 ;
  RECT 46.280 178.640 49.820 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 32.640 178.640 36.180 179.760 ;
  LAYER metal4 ;
  RECT 32.640 178.640 36.180 179.760 ;
  LAYER metal3 ;
  RECT 32.640 178.640 36.180 179.760 ;
  LAYER metal2 ;
  RECT 32.640 178.640 36.180 179.760 ;
  LAYER metal1 ;
  RECT 32.640 178.640 36.180 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 21.480 178.640 25.020 179.760 ;
  LAYER metal4 ;
  RECT 21.480 178.640 25.020 179.760 ;
  LAYER metal3 ;
  RECT 21.480 178.640 25.020 179.760 ;
  LAYER metal2 ;
  RECT 21.480 178.640 25.020 179.760 ;
  LAYER metal1 ;
  RECT 21.480 178.640 25.020 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 7.220 178.640 10.760 179.760 ;
  LAYER metal4 ;
  RECT 7.220 178.640 10.760 179.760 ;
  LAYER metal3 ;
  RECT 7.220 178.640 10.760 179.760 ;
  LAYER metal2 ;
  RECT 7.220 178.640 10.760 179.760 ;
  LAYER metal1 ;
  RECT 7.220 178.640 10.760 179.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3535.640 0.000 3539.180 1.120 ;
  LAYER metal4 ;
  RECT 3535.640 0.000 3539.180 1.120 ;
  LAYER metal3 ;
  RECT 3535.640 0.000 3539.180 1.120 ;
  LAYER metal2 ;
  RECT 3535.640 0.000 3539.180 1.120 ;
  LAYER metal1 ;
  RECT 3535.640 0.000 3539.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3526.960 0.000 3530.500 1.120 ;
  LAYER metal4 ;
  RECT 3526.960 0.000 3530.500 1.120 ;
  LAYER metal3 ;
  RECT 3526.960 0.000 3530.500 1.120 ;
  LAYER metal2 ;
  RECT 3526.960 0.000 3530.500 1.120 ;
  LAYER metal1 ;
  RECT 3526.960 0.000 3530.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3513.320 0.000 3516.860 1.120 ;
  LAYER metal4 ;
  RECT 3513.320 0.000 3516.860 1.120 ;
  LAYER metal3 ;
  RECT 3513.320 0.000 3516.860 1.120 ;
  LAYER metal2 ;
  RECT 3513.320 0.000 3516.860 1.120 ;
  LAYER metal1 ;
  RECT 3513.320 0.000 3516.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3446.360 0.000 3449.900 1.120 ;
  LAYER metal4 ;
  RECT 3446.360 0.000 3449.900 1.120 ;
  LAYER metal3 ;
  RECT 3446.360 0.000 3449.900 1.120 ;
  LAYER metal2 ;
  RECT 3446.360 0.000 3449.900 1.120 ;
  LAYER metal1 ;
  RECT 3446.360 0.000 3449.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3432.720 0.000 3436.260 1.120 ;
  LAYER metal4 ;
  RECT 3432.720 0.000 3436.260 1.120 ;
  LAYER metal3 ;
  RECT 3432.720 0.000 3436.260 1.120 ;
  LAYER metal2 ;
  RECT 3432.720 0.000 3436.260 1.120 ;
  LAYER metal1 ;
  RECT 3432.720 0.000 3436.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3419.080 0.000 3422.620 1.120 ;
  LAYER metal4 ;
  RECT 3419.080 0.000 3422.620 1.120 ;
  LAYER metal3 ;
  RECT 3419.080 0.000 3422.620 1.120 ;
  LAYER metal2 ;
  RECT 3419.080 0.000 3422.620 1.120 ;
  LAYER metal1 ;
  RECT 3419.080 0.000 3422.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3406.060 0.000 3409.600 1.120 ;
  LAYER metal4 ;
  RECT 3406.060 0.000 3409.600 1.120 ;
  LAYER metal3 ;
  RECT 3406.060 0.000 3409.600 1.120 ;
  LAYER metal2 ;
  RECT 3406.060 0.000 3409.600 1.120 ;
  LAYER metal1 ;
  RECT 3406.060 0.000 3409.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3392.420 0.000 3395.960 1.120 ;
  LAYER metal4 ;
  RECT 3392.420 0.000 3395.960 1.120 ;
  LAYER metal3 ;
  RECT 3392.420 0.000 3395.960 1.120 ;
  LAYER metal2 ;
  RECT 3392.420 0.000 3395.960 1.120 ;
  LAYER metal1 ;
  RECT 3392.420 0.000 3395.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3378.780 0.000 3382.320 1.120 ;
  LAYER metal4 ;
  RECT 3378.780 0.000 3382.320 1.120 ;
  LAYER metal3 ;
  RECT 3378.780 0.000 3382.320 1.120 ;
  LAYER metal2 ;
  RECT 3378.780 0.000 3382.320 1.120 ;
  LAYER metal1 ;
  RECT 3378.780 0.000 3382.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3311.820 0.000 3315.360 1.120 ;
  LAYER metal4 ;
  RECT 3311.820 0.000 3315.360 1.120 ;
  LAYER metal3 ;
  RECT 3311.820 0.000 3315.360 1.120 ;
  LAYER metal2 ;
  RECT 3311.820 0.000 3315.360 1.120 ;
  LAYER metal1 ;
  RECT 3311.820 0.000 3315.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3298.180 0.000 3301.720 1.120 ;
  LAYER metal4 ;
  RECT 3298.180 0.000 3301.720 1.120 ;
  LAYER metal3 ;
  RECT 3298.180 0.000 3301.720 1.120 ;
  LAYER metal2 ;
  RECT 3298.180 0.000 3301.720 1.120 ;
  LAYER metal1 ;
  RECT 3298.180 0.000 3301.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3284.540 0.000 3288.080 1.120 ;
  LAYER metal4 ;
  RECT 3284.540 0.000 3288.080 1.120 ;
  LAYER metal3 ;
  RECT 3284.540 0.000 3288.080 1.120 ;
  LAYER metal2 ;
  RECT 3284.540 0.000 3288.080 1.120 ;
  LAYER metal1 ;
  RECT 3284.540 0.000 3288.080 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3271.520 0.000 3275.060 1.120 ;
  LAYER metal4 ;
  RECT 3271.520 0.000 3275.060 1.120 ;
  LAYER metal3 ;
  RECT 3271.520 0.000 3275.060 1.120 ;
  LAYER metal2 ;
  RECT 3271.520 0.000 3275.060 1.120 ;
  LAYER metal1 ;
  RECT 3271.520 0.000 3275.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3257.880 0.000 3261.420 1.120 ;
  LAYER metal4 ;
  RECT 3257.880 0.000 3261.420 1.120 ;
  LAYER metal3 ;
  RECT 3257.880 0.000 3261.420 1.120 ;
  LAYER metal2 ;
  RECT 3257.880 0.000 3261.420 1.120 ;
  LAYER metal1 ;
  RECT 3257.880 0.000 3261.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3244.240 0.000 3247.780 1.120 ;
  LAYER metal4 ;
  RECT 3244.240 0.000 3247.780 1.120 ;
  LAYER metal3 ;
  RECT 3244.240 0.000 3247.780 1.120 ;
  LAYER metal2 ;
  RECT 3244.240 0.000 3247.780 1.120 ;
  LAYER metal1 ;
  RECT 3244.240 0.000 3247.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3177.280 0.000 3180.820 1.120 ;
  LAYER metal4 ;
  RECT 3177.280 0.000 3180.820 1.120 ;
  LAYER metal3 ;
  RECT 3177.280 0.000 3180.820 1.120 ;
  LAYER metal2 ;
  RECT 3177.280 0.000 3180.820 1.120 ;
  LAYER metal1 ;
  RECT 3177.280 0.000 3180.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3163.640 0.000 3167.180 1.120 ;
  LAYER metal4 ;
  RECT 3163.640 0.000 3167.180 1.120 ;
  LAYER metal3 ;
  RECT 3163.640 0.000 3167.180 1.120 ;
  LAYER metal2 ;
  RECT 3163.640 0.000 3167.180 1.120 ;
  LAYER metal1 ;
  RECT 3163.640 0.000 3167.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3150.620 0.000 3154.160 1.120 ;
  LAYER metal4 ;
  RECT 3150.620 0.000 3154.160 1.120 ;
  LAYER metal3 ;
  RECT 3150.620 0.000 3154.160 1.120 ;
  LAYER metal2 ;
  RECT 3150.620 0.000 3154.160 1.120 ;
  LAYER metal1 ;
  RECT 3150.620 0.000 3154.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3136.980 0.000 3140.520 1.120 ;
  LAYER metal4 ;
  RECT 3136.980 0.000 3140.520 1.120 ;
  LAYER metal3 ;
  RECT 3136.980 0.000 3140.520 1.120 ;
  LAYER metal2 ;
  RECT 3136.980 0.000 3140.520 1.120 ;
  LAYER metal1 ;
  RECT 3136.980 0.000 3140.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3123.340 0.000 3126.880 1.120 ;
  LAYER metal4 ;
  RECT 3123.340 0.000 3126.880 1.120 ;
  LAYER metal3 ;
  RECT 3123.340 0.000 3126.880 1.120 ;
  LAYER metal2 ;
  RECT 3123.340 0.000 3126.880 1.120 ;
  LAYER metal1 ;
  RECT 3123.340 0.000 3126.880 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3112.180 0.000 3115.720 1.120 ;
  LAYER metal4 ;
  RECT 3112.180 0.000 3115.720 1.120 ;
  LAYER metal3 ;
  RECT 3112.180 0.000 3115.720 1.120 ;
  LAYER metal2 ;
  RECT 3112.180 0.000 3115.720 1.120 ;
  LAYER metal1 ;
  RECT 3112.180 0.000 3115.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3042.740 0.000 3046.280 1.120 ;
  LAYER metal4 ;
  RECT 3042.740 0.000 3046.280 1.120 ;
  LAYER metal3 ;
  RECT 3042.740 0.000 3046.280 1.120 ;
  LAYER metal2 ;
  RECT 3042.740 0.000 3046.280 1.120 ;
  LAYER metal1 ;
  RECT 3042.740 0.000 3046.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3029.720 0.000 3033.260 1.120 ;
  LAYER metal4 ;
  RECT 3029.720 0.000 3033.260 1.120 ;
  LAYER metal3 ;
  RECT 3029.720 0.000 3033.260 1.120 ;
  LAYER metal2 ;
  RECT 3029.720 0.000 3033.260 1.120 ;
  LAYER metal1 ;
  RECT 3029.720 0.000 3033.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3016.080 0.000 3019.620 1.120 ;
  LAYER metal4 ;
  RECT 3016.080 0.000 3019.620 1.120 ;
  LAYER metal3 ;
  RECT 3016.080 0.000 3019.620 1.120 ;
  LAYER metal2 ;
  RECT 3016.080 0.000 3019.620 1.120 ;
  LAYER metal1 ;
  RECT 3016.080 0.000 3019.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3002.440 0.000 3005.980 1.120 ;
  LAYER metal4 ;
  RECT 3002.440 0.000 3005.980 1.120 ;
  LAYER metal3 ;
  RECT 3002.440 0.000 3005.980 1.120 ;
  LAYER metal2 ;
  RECT 3002.440 0.000 3005.980 1.120 ;
  LAYER metal1 ;
  RECT 3002.440 0.000 3005.980 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2989.420 0.000 2992.960 1.120 ;
  LAYER metal4 ;
  RECT 2989.420 0.000 2992.960 1.120 ;
  LAYER metal3 ;
  RECT 2989.420 0.000 2992.960 1.120 ;
  LAYER metal2 ;
  RECT 2989.420 0.000 2992.960 1.120 ;
  LAYER metal1 ;
  RECT 2989.420 0.000 2992.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2975.780 0.000 2979.320 1.120 ;
  LAYER metal4 ;
  RECT 2975.780 0.000 2979.320 1.120 ;
  LAYER metal3 ;
  RECT 2975.780 0.000 2979.320 1.120 ;
  LAYER metal2 ;
  RECT 2975.780 0.000 2979.320 1.120 ;
  LAYER metal1 ;
  RECT 2975.780 0.000 2979.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2908.200 0.000 2911.740 1.120 ;
  LAYER metal4 ;
  RECT 2908.200 0.000 2911.740 1.120 ;
  LAYER metal3 ;
  RECT 2908.200 0.000 2911.740 1.120 ;
  LAYER metal2 ;
  RECT 2908.200 0.000 2911.740 1.120 ;
  LAYER metal1 ;
  RECT 2908.200 0.000 2911.740 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2895.180 0.000 2898.720 1.120 ;
  LAYER metal4 ;
  RECT 2895.180 0.000 2898.720 1.120 ;
  LAYER metal3 ;
  RECT 2895.180 0.000 2898.720 1.120 ;
  LAYER metal2 ;
  RECT 2895.180 0.000 2898.720 1.120 ;
  LAYER metal1 ;
  RECT 2895.180 0.000 2898.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2881.540 0.000 2885.080 1.120 ;
  LAYER metal4 ;
  RECT 2881.540 0.000 2885.080 1.120 ;
  LAYER metal3 ;
  RECT 2881.540 0.000 2885.080 1.120 ;
  LAYER metal2 ;
  RECT 2881.540 0.000 2885.080 1.120 ;
  LAYER metal1 ;
  RECT 2881.540 0.000 2885.080 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2867.900 0.000 2871.440 1.120 ;
  LAYER metal4 ;
  RECT 2867.900 0.000 2871.440 1.120 ;
  LAYER metal3 ;
  RECT 2867.900 0.000 2871.440 1.120 ;
  LAYER metal2 ;
  RECT 2867.900 0.000 2871.440 1.120 ;
  LAYER metal1 ;
  RECT 2867.900 0.000 2871.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2854.880 0.000 2858.420 1.120 ;
  LAYER metal4 ;
  RECT 2854.880 0.000 2858.420 1.120 ;
  LAYER metal3 ;
  RECT 2854.880 0.000 2858.420 1.120 ;
  LAYER metal2 ;
  RECT 2854.880 0.000 2858.420 1.120 ;
  LAYER metal1 ;
  RECT 2854.880 0.000 2858.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2841.240 0.000 2844.780 1.120 ;
  LAYER metal4 ;
  RECT 2841.240 0.000 2844.780 1.120 ;
  LAYER metal3 ;
  RECT 2841.240 0.000 2844.780 1.120 ;
  LAYER metal2 ;
  RECT 2841.240 0.000 2844.780 1.120 ;
  LAYER metal1 ;
  RECT 2841.240 0.000 2844.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2774.280 0.000 2777.820 1.120 ;
  LAYER metal4 ;
  RECT 2774.280 0.000 2777.820 1.120 ;
  LAYER metal3 ;
  RECT 2774.280 0.000 2777.820 1.120 ;
  LAYER metal2 ;
  RECT 2774.280 0.000 2777.820 1.120 ;
  LAYER metal1 ;
  RECT 2774.280 0.000 2777.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2760.640 0.000 2764.180 1.120 ;
  LAYER metal4 ;
  RECT 2760.640 0.000 2764.180 1.120 ;
  LAYER metal3 ;
  RECT 2760.640 0.000 2764.180 1.120 ;
  LAYER metal2 ;
  RECT 2760.640 0.000 2764.180 1.120 ;
  LAYER metal1 ;
  RECT 2760.640 0.000 2764.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2747.000 0.000 2750.540 1.120 ;
  LAYER metal4 ;
  RECT 2747.000 0.000 2750.540 1.120 ;
  LAYER metal3 ;
  RECT 2747.000 0.000 2750.540 1.120 ;
  LAYER metal2 ;
  RECT 2747.000 0.000 2750.540 1.120 ;
  LAYER metal1 ;
  RECT 2747.000 0.000 2750.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2733.980 0.000 2737.520 1.120 ;
  LAYER metal4 ;
  RECT 2733.980 0.000 2737.520 1.120 ;
  LAYER metal3 ;
  RECT 2733.980 0.000 2737.520 1.120 ;
  LAYER metal2 ;
  RECT 2733.980 0.000 2737.520 1.120 ;
  LAYER metal1 ;
  RECT 2733.980 0.000 2737.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2720.340 0.000 2723.880 1.120 ;
  LAYER metal4 ;
  RECT 2720.340 0.000 2723.880 1.120 ;
  LAYER metal3 ;
  RECT 2720.340 0.000 2723.880 1.120 ;
  LAYER metal2 ;
  RECT 2720.340 0.000 2723.880 1.120 ;
  LAYER metal1 ;
  RECT 2720.340 0.000 2723.880 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2706.700 0.000 2710.240 1.120 ;
  LAYER metal4 ;
  RECT 2706.700 0.000 2710.240 1.120 ;
  LAYER metal3 ;
  RECT 2706.700 0.000 2710.240 1.120 ;
  LAYER metal2 ;
  RECT 2706.700 0.000 2710.240 1.120 ;
  LAYER metal1 ;
  RECT 2706.700 0.000 2710.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2639.740 0.000 2643.280 1.120 ;
  LAYER metal4 ;
  RECT 2639.740 0.000 2643.280 1.120 ;
  LAYER metal3 ;
  RECT 2639.740 0.000 2643.280 1.120 ;
  LAYER metal2 ;
  RECT 2639.740 0.000 2643.280 1.120 ;
  LAYER metal1 ;
  RECT 2639.740 0.000 2643.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2626.100 0.000 2629.640 1.120 ;
  LAYER metal4 ;
  RECT 2626.100 0.000 2629.640 1.120 ;
  LAYER metal3 ;
  RECT 2626.100 0.000 2629.640 1.120 ;
  LAYER metal2 ;
  RECT 2626.100 0.000 2629.640 1.120 ;
  LAYER metal1 ;
  RECT 2626.100 0.000 2629.640 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2613.080 0.000 2616.620 1.120 ;
  LAYER metal4 ;
  RECT 2613.080 0.000 2616.620 1.120 ;
  LAYER metal3 ;
  RECT 2613.080 0.000 2616.620 1.120 ;
  LAYER metal2 ;
  RECT 2613.080 0.000 2616.620 1.120 ;
  LAYER metal1 ;
  RECT 2613.080 0.000 2616.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2599.440 0.000 2602.980 1.120 ;
  LAYER metal4 ;
  RECT 2599.440 0.000 2602.980 1.120 ;
  LAYER metal3 ;
  RECT 2599.440 0.000 2602.980 1.120 ;
  LAYER metal2 ;
  RECT 2599.440 0.000 2602.980 1.120 ;
  LAYER metal1 ;
  RECT 2599.440 0.000 2602.980 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2585.800 0.000 2589.340 1.120 ;
  LAYER metal4 ;
  RECT 2585.800 0.000 2589.340 1.120 ;
  LAYER metal3 ;
  RECT 2585.800 0.000 2589.340 1.120 ;
  LAYER metal2 ;
  RECT 2585.800 0.000 2589.340 1.120 ;
  LAYER metal1 ;
  RECT 2585.800 0.000 2589.340 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2572.780 0.000 2576.320 1.120 ;
  LAYER metal4 ;
  RECT 2572.780 0.000 2576.320 1.120 ;
  LAYER metal3 ;
  RECT 2572.780 0.000 2576.320 1.120 ;
  LAYER metal2 ;
  RECT 2572.780 0.000 2576.320 1.120 ;
  LAYER metal1 ;
  RECT 2572.780 0.000 2576.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2505.200 0.000 2508.740 1.120 ;
  LAYER metal4 ;
  RECT 2505.200 0.000 2508.740 1.120 ;
  LAYER metal3 ;
  RECT 2505.200 0.000 2508.740 1.120 ;
  LAYER metal2 ;
  RECT 2505.200 0.000 2508.740 1.120 ;
  LAYER metal1 ;
  RECT 2505.200 0.000 2508.740 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2491.560 0.000 2495.100 1.120 ;
  LAYER metal4 ;
  RECT 2491.560 0.000 2495.100 1.120 ;
  LAYER metal3 ;
  RECT 2491.560 0.000 2495.100 1.120 ;
  LAYER metal2 ;
  RECT 2491.560 0.000 2495.100 1.120 ;
  LAYER metal1 ;
  RECT 2491.560 0.000 2495.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2478.540 0.000 2482.080 1.120 ;
  LAYER metal4 ;
  RECT 2478.540 0.000 2482.080 1.120 ;
  LAYER metal3 ;
  RECT 2478.540 0.000 2482.080 1.120 ;
  LAYER metal2 ;
  RECT 2478.540 0.000 2482.080 1.120 ;
  LAYER metal1 ;
  RECT 2478.540 0.000 2482.080 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2464.900 0.000 2468.440 1.120 ;
  LAYER metal4 ;
  RECT 2464.900 0.000 2468.440 1.120 ;
  LAYER metal3 ;
  RECT 2464.900 0.000 2468.440 1.120 ;
  LAYER metal2 ;
  RECT 2464.900 0.000 2468.440 1.120 ;
  LAYER metal1 ;
  RECT 2464.900 0.000 2468.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2451.260 0.000 2454.800 1.120 ;
  LAYER metal4 ;
  RECT 2451.260 0.000 2454.800 1.120 ;
  LAYER metal3 ;
  RECT 2451.260 0.000 2454.800 1.120 ;
  LAYER metal2 ;
  RECT 2451.260 0.000 2454.800 1.120 ;
  LAYER metal1 ;
  RECT 2451.260 0.000 2454.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2438.240 0.000 2441.780 1.120 ;
  LAYER metal4 ;
  RECT 2438.240 0.000 2441.780 1.120 ;
  LAYER metal3 ;
  RECT 2438.240 0.000 2441.780 1.120 ;
  LAYER metal2 ;
  RECT 2438.240 0.000 2441.780 1.120 ;
  LAYER metal1 ;
  RECT 2438.240 0.000 2441.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2370.660 0.000 2374.200 1.120 ;
  LAYER metal4 ;
  RECT 2370.660 0.000 2374.200 1.120 ;
  LAYER metal3 ;
  RECT 2370.660 0.000 2374.200 1.120 ;
  LAYER metal2 ;
  RECT 2370.660 0.000 2374.200 1.120 ;
  LAYER metal1 ;
  RECT 2370.660 0.000 2374.200 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2357.640 0.000 2361.180 1.120 ;
  LAYER metal4 ;
  RECT 2357.640 0.000 2361.180 1.120 ;
  LAYER metal3 ;
  RECT 2357.640 0.000 2361.180 1.120 ;
  LAYER metal2 ;
  RECT 2357.640 0.000 2361.180 1.120 ;
  LAYER metal1 ;
  RECT 2357.640 0.000 2361.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2344.000 0.000 2347.540 1.120 ;
  LAYER metal4 ;
  RECT 2344.000 0.000 2347.540 1.120 ;
  LAYER metal3 ;
  RECT 2344.000 0.000 2347.540 1.120 ;
  LAYER metal2 ;
  RECT 2344.000 0.000 2347.540 1.120 ;
  LAYER metal1 ;
  RECT 2344.000 0.000 2347.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2330.360 0.000 2333.900 1.120 ;
  LAYER metal4 ;
  RECT 2330.360 0.000 2333.900 1.120 ;
  LAYER metal3 ;
  RECT 2330.360 0.000 2333.900 1.120 ;
  LAYER metal2 ;
  RECT 2330.360 0.000 2333.900 1.120 ;
  LAYER metal1 ;
  RECT 2330.360 0.000 2333.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2317.340 0.000 2320.880 1.120 ;
  LAYER metal4 ;
  RECT 2317.340 0.000 2320.880 1.120 ;
  LAYER metal3 ;
  RECT 2317.340 0.000 2320.880 1.120 ;
  LAYER metal2 ;
  RECT 2317.340 0.000 2320.880 1.120 ;
  LAYER metal1 ;
  RECT 2317.340 0.000 2320.880 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2303.700 0.000 2307.240 1.120 ;
  LAYER metal4 ;
  RECT 2303.700 0.000 2307.240 1.120 ;
  LAYER metal3 ;
  RECT 2303.700 0.000 2307.240 1.120 ;
  LAYER metal2 ;
  RECT 2303.700 0.000 2307.240 1.120 ;
  LAYER metal1 ;
  RECT 2303.700 0.000 2307.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2236.740 0.000 2240.280 1.120 ;
  LAYER metal4 ;
  RECT 2236.740 0.000 2240.280 1.120 ;
  LAYER metal3 ;
  RECT 2236.740 0.000 2240.280 1.120 ;
  LAYER metal2 ;
  RECT 2236.740 0.000 2240.280 1.120 ;
  LAYER metal1 ;
  RECT 2236.740 0.000 2240.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2223.100 0.000 2226.640 1.120 ;
  LAYER metal4 ;
  RECT 2223.100 0.000 2226.640 1.120 ;
  LAYER metal3 ;
  RECT 2223.100 0.000 2226.640 1.120 ;
  LAYER metal2 ;
  RECT 2223.100 0.000 2226.640 1.120 ;
  LAYER metal1 ;
  RECT 2223.100 0.000 2226.640 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2209.460 0.000 2213.000 1.120 ;
  LAYER metal4 ;
  RECT 2209.460 0.000 2213.000 1.120 ;
  LAYER metal3 ;
  RECT 2209.460 0.000 2213.000 1.120 ;
  LAYER metal2 ;
  RECT 2209.460 0.000 2213.000 1.120 ;
  LAYER metal1 ;
  RECT 2209.460 0.000 2213.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2196.440 0.000 2199.980 1.120 ;
  LAYER metal4 ;
  RECT 2196.440 0.000 2199.980 1.120 ;
  LAYER metal3 ;
  RECT 2196.440 0.000 2199.980 1.120 ;
  LAYER metal2 ;
  RECT 2196.440 0.000 2199.980 1.120 ;
  LAYER metal1 ;
  RECT 2196.440 0.000 2199.980 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2182.800 0.000 2186.340 1.120 ;
  LAYER metal4 ;
  RECT 2182.800 0.000 2186.340 1.120 ;
  LAYER metal3 ;
  RECT 2182.800 0.000 2186.340 1.120 ;
  LAYER metal2 ;
  RECT 2182.800 0.000 2186.340 1.120 ;
  LAYER metal1 ;
  RECT 2182.800 0.000 2186.340 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2169.160 0.000 2172.700 1.120 ;
  LAYER metal4 ;
  RECT 2169.160 0.000 2172.700 1.120 ;
  LAYER metal3 ;
  RECT 2169.160 0.000 2172.700 1.120 ;
  LAYER metal2 ;
  RECT 2169.160 0.000 2172.700 1.120 ;
  LAYER metal1 ;
  RECT 2169.160 0.000 2172.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2102.200 0.000 2105.740 1.120 ;
  LAYER metal4 ;
  RECT 2102.200 0.000 2105.740 1.120 ;
  LAYER metal3 ;
  RECT 2102.200 0.000 2105.740 1.120 ;
  LAYER metal2 ;
  RECT 2102.200 0.000 2105.740 1.120 ;
  LAYER metal1 ;
  RECT 2102.200 0.000 2105.740 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2088.560 0.000 2092.100 1.120 ;
  LAYER metal4 ;
  RECT 2088.560 0.000 2092.100 1.120 ;
  LAYER metal3 ;
  RECT 2088.560 0.000 2092.100 1.120 ;
  LAYER metal2 ;
  RECT 2088.560 0.000 2092.100 1.120 ;
  LAYER metal1 ;
  RECT 2088.560 0.000 2092.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2074.920 0.000 2078.460 1.120 ;
  LAYER metal4 ;
  RECT 2074.920 0.000 2078.460 1.120 ;
  LAYER metal3 ;
  RECT 2074.920 0.000 2078.460 1.120 ;
  LAYER metal2 ;
  RECT 2074.920 0.000 2078.460 1.120 ;
  LAYER metal1 ;
  RECT 2074.920 0.000 2078.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2061.900 0.000 2065.440 1.120 ;
  LAYER metal4 ;
  RECT 2061.900 0.000 2065.440 1.120 ;
  LAYER metal3 ;
  RECT 2061.900 0.000 2065.440 1.120 ;
  LAYER metal2 ;
  RECT 2061.900 0.000 2065.440 1.120 ;
  LAYER metal1 ;
  RECT 2061.900 0.000 2065.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2048.260 0.000 2051.800 1.120 ;
  LAYER metal4 ;
  RECT 2048.260 0.000 2051.800 1.120 ;
  LAYER metal3 ;
  RECT 2048.260 0.000 2051.800 1.120 ;
  LAYER metal2 ;
  RECT 2048.260 0.000 2051.800 1.120 ;
  LAYER metal1 ;
  RECT 2048.260 0.000 2051.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2034.620 0.000 2038.160 1.120 ;
  LAYER metal4 ;
  RECT 2034.620 0.000 2038.160 1.120 ;
  LAYER metal3 ;
  RECT 2034.620 0.000 2038.160 1.120 ;
  LAYER metal2 ;
  RECT 2034.620 0.000 2038.160 1.120 ;
  LAYER metal1 ;
  RECT 2034.620 0.000 2038.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1967.660 0.000 1971.200 1.120 ;
  LAYER metal4 ;
  RECT 1967.660 0.000 1971.200 1.120 ;
  LAYER metal3 ;
  RECT 1967.660 0.000 1971.200 1.120 ;
  LAYER metal2 ;
  RECT 1967.660 0.000 1971.200 1.120 ;
  LAYER metal1 ;
  RECT 1967.660 0.000 1971.200 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1954.020 0.000 1957.560 1.120 ;
  LAYER metal4 ;
  RECT 1954.020 0.000 1957.560 1.120 ;
  LAYER metal3 ;
  RECT 1954.020 0.000 1957.560 1.120 ;
  LAYER metal2 ;
  RECT 1954.020 0.000 1957.560 1.120 ;
  LAYER metal1 ;
  RECT 1954.020 0.000 1957.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1941.000 0.000 1944.540 1.120 ;
  LAYER metal4 ;
  RECT 1941.000 0.000 1944.540 1.120 ;
  LAYER metal3 ;
  RECT 1941.000 0.000 1944.540 1.120 ;
  LAYER metal2 ;
  RECT 1941.000 0.000 1944.540 1.120 ;
  LAYER metal1 ;
  RECT 1941.000 0.000 1944.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1927.360 0.000 1930.900 1.120 ;
  LAYER metal4 ;
  RECT 1927.360 0.000 1930.900 1.120 ;
  LAYER metal3 ;
  RECT 1927.360 0.000 1930.900 1.120 ;
  LAYER metal2 ;
  RECT 1927.360 0.000 1930.900 1.120 ;
  LAYER metal1 ;
  RECT 1927.360 0.000 1930.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1913.720 0.000 1917.260 1.120 ;
  LAYER metal4 ;
  RECT 1913.720 0.000 1917.260 1.120 ;
  LAYER metal3 ;
  RECT 1913.720 0.000 1917.260 1.120 ;
  LAYER metal2 ;
  RECT 1913.720 0.000 1917.260 1.120 ;
  LAYER metal1 ;
  RECT 1913.720 0.000 1917.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1900.700 0.000 1904.240 1.120 ;
  LAYER metal4 ;
  RECT 1900.700 0.000 1904.240 1.120 ;
  LAYER metal3 ;
  RECT 1900.700 0.000 1904.240 1.120 ;
  LAYER metal2 ;
  RECT 1900.700 0.000 1904.240 1.120 ;
  LAYER metal1 ;
  RECT 1900.700 0.000 1904.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1833.120 0.000 1836.660 1.120 ;
  LAYER metal4 ;
  RECT 1833.120 0.000 1836.660 1.120 ;
  LAYER metal3 ;
  RECT 1833.120 0.000 1836.660 1.120 ;
  LAYER metal2 ;
  RECT 1833.120 0.000 1836.660 1.120 ;
  LAYER metal1 ;
  RECT 1833.120 0.000 1836.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1821.960 0.000 1825.500 1.120 ;
  LAYER metal4 ;
  RECT 1821.960 0.000 1825.500 1.120 ;
  LAYER metal3 ;
  RECT 1821.960 0.000 1825.500 1.120 ;
  LAYER metal2 ;
  RECT 1821.960 0.000 1825.500 1.120 ;
  LAYER metal1 ;
  RECT 1821.960 0.000 1825.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1805.840 0.000 1809.380 1.120 ;
  LAYER metal4 ;
  RECT 1805.840 0.000 1809.380 1.120 ;
  LAYER metal3 ;
  RECT 1805.840 0.000 1809.380 1.120 ;
  LAYER metal2 ;
  RECT 1805.840 0.000 1809.380 1.120 ;
  LAYER metal1 ;
  RECT 1805.840 0.000 1809.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1797.160 0.000 1800.700 1.120 ;
  LAYER metal4 ;
  RECT 1797.160 0.000 1800.700 1.120 ;
  LAYER metal3 ;
  RECT 1797.160 0.000 1800.700 1.120 ;
  LAYER metal2 ;
  RECT 1797.160 0.000 1800.700 1.120 ;
  LAYER metal1 ;
  RECT 1797.160 0.000 1800.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1784.140 0.000 1787.680 1.120 ;
  LAYER metal4 ;
  RECT 1784.140 0.000 1787.680 1.120 ;
  LAYER metal3 ;
  RECT 1784.140 0.000 1787.680 1.120 ;
  LAYER metal2 ;
  RECT 1784.140 0.000 1787.680 1.120 ;
  LAYER metal1 ;
  RECT 1784.140 0.000 1787.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1771.120 0.000 1774.660 1.120 ;
  LAYER metal4 ;
  RECT 1771.120 0.000 1774.660 1.120 ;
  LAYER metal3 ;
  RECT 1771.120 0.000 1774.660 1.120 ;
  LAYER metal2 ;
  RECT 1771.120 0.000 1774.660 1.120 ;
  LAYER metal1 ;
  RECT 1771.120 0.000 1774.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1685.560 0.000 1689.100 1.120 ;
  LAYER metal4 ;
  RECT 1685.560 0.000 1689.100 1.120 ;
  LAYER metal3 ;
  RECT 1685.560 0.000 1689.100 1.120 ;
  LAYER metal2 ;
  RECT 1685.560 0.000 1689.100 1.120 ;
  LAYER metal1 ;
  RECT 1685.560 0.000 1689.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1672.540 0.000 1676.080 1.120 ;
  LAYER metal4 ;
  RECT 1672.540 0.000 1676.080 1.120 ;
  LAYER metal3 ;
  RECT 1672.540 0.000 1676.080 1.120 ;
  LAYER metal2 ;
  RECT 1672.540 0.000 1676.080 1.120 ;
  LAYER metal1 ;
  RECT 1672.540 0.000 1676.080 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1658.900 0.000 1662.440 1.120 ;
  LAYER metal4 ;
  RECT 1658.900 0.000 1662.440 1.120 ;
  LAYER metal3 ;
  RECT 1658.900 0.000 1662.440 1.120 ;
  LAYER metal2 ;
  RECT 1658.900 0.000 1662.440 1.120 ;
  LAYER metal1 ;
  RECT 1658.900 0.000 1662.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1645.260 0.000 1648.800 1.120 ;
  LAYER metal4 ;
  RECT 1645.260 0.000 1648.800 1.120 ;
  LAYER metal3 ;
  RECT 1645.260 0.000 1648.800 1.120 ;
  LAYER metal2 ;
  RECT 1645.260 0.000 1648.800 1.120 ;
  LAYER metal1 ;
  RECT 1645.260 0.000 1648.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1632.240 0.000 1635.780 1.120 ;
  LAYER metal4 ;
  RECT 1632.240 0.000 1635.780 1.120 ;
  LAYER metal3 ;
  RECT 1632.240 0.000 1635.780 1.120 ;
  LAYER metal2 ;
  RECT 1632.240 0.000 1635.780 1.120 ;
  LAYER metal1 ;
  RECT 1632.240 0.000 1635.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1618.600 0.000 1622.140 1.120 ;
  LAYER metal4 ;
  RECT 1618.600 0.000 1622.140 1.120 ;
  LAYER metal3 ;
  RECT 1618.600 0.000 1622.140 1.120 ;
  LAYER metal2 ;
  RECT 1618.600 0.000 1622.140 1.120 ;
  LAYER metal1 ;
  RECT 1618.600 0.000 1622.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1551.640 0.000 1555.180 1.120 ;
  LAYER metal4 ;
  RECT 1551.640 0.000 1555.180 1.120 ;
  LAYER metal3 ;
  RECT 1551.640 0.000 1555.180 1.120 ;
  LAYER metal2 ;
  RECT 1551.640 0.000 1555.180 1.120 ;
  LAYER metal1 ;
  RECT 1551.640 0.000 1555.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1538.000 0.000 1541.540 1.120 ;
  LAYER metal4 ;
  RECT 1538.000 0.000 1541.540 1.120 ;
  LAYER metal3 ;
  RECT 1538.000 0.000 1541.540 1.120 ;
  LAYER metal2 ;
  RECT 1538.000 0.000 1541.540 1.120 ;
  LAYER metal1 ;
  RECT 1538.000 0.000 1541.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1524.360 0.000 1527.900 1.120 ;
  LAYER metal4 ;
  RECT 1524.360 0.000 1527.900 1.120 ;
  LAYER metal3 ;
  RECT 1524.360 0.000 1527.900 1.120 ;
  LAYER metal2 ;
  RECT 1524.360 0.000 1527.900 1.120 ;
  LAYER metal1 ;
  RECT 1524.360 0.000 1527.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1511.340 0.000 1514.880 1.120 ;
  LAYER metal4 ;
  RECT 1511.340 0.000 1514.880 1.120 ;
  LAYER metal3 ;
  RECT 1511.340 0.000 1514.880 1.120 ;
  LAYER metal2 ;
  RECT 1511.340 0.000 1514.880 1.120 ;
  LAYER metal1 ;
  RECT 1511.340 0.000 1514.880 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1497.700 0.000 1501.240 1.120 ;
  LAYER metal4 ;
  RECT 1497.700 0.000 1501.240 1.120 ;
  LAYER metal3 ;
  RECT 1497.700 0.000 1501.240 1.120 ;
  LAYER metal2 ;
  RECT 1497.700 0.000 1501.240 1.120 ;
  LAYER metal1 ;
  RECT 1497.700 0.000 1501.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1484.060 0.000 1487.600 1.120 ;
  LAYER metal4 ;
  RECT 1484.060 0.000 1487.600 1.120 ;
  LAYER metal3 ;
  RECT 1484.060 0.000 1487.600 1.120 ;
  LAYER metal2 ;
  RECT 1484.060 0.000 1487.600 1.120 ;
  LAYER metal1 ;
  RECT 1484.060 0.000 1487.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1417.100 0.000 1420.640 1.120 ;
  LAYER metal4 ;
  RECT 1417.100 0.000 1420.640 1.120 ;
  LAYER metal3 ;
  RECT 1417.100 0.000 1420.640 1.120 ;
  LAYER metal2 ;
  RECT 1417.100 0.000 1420.640 1.120 ;
  LAYER metal1 ;
  RECT 1417.100 0.000 1420.640 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1403.460 0.000 1407.000 1.120 ;
  LAYER metal4 ;
  RECT 1403.460 0.000 1407.000 1.120 ;
  LAYER metal3 ;
  RECT 1403.460 0.000 1407.000 1.120 ;
  LAYER metal2 ;
  RECT 1403.460 0.000 1407.000 1.120 ;
  LAYER metal1 ;
  RECT 1403.460 0.000 1407.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1390.440 0.000 1393.980 1.120 ;
  LAYER metal4 ;
  RECT 1390.440 0.000 1393.980 1.120 ;
  LAYER metal3 ;
  RECT 1390.440 0.000 1393.980 1.120 ;
  LAYER metal2 ;
  RECT 1390.440 0.000 1393.980 1.120 ;
  LAYER metal1 ;
  RECT 1390.440 0.000 1393.980 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1376.800 0.000 1380.340 1.120 ;
  LAYER metal4 ;
  RECT 1376.800 0.000 1380.340 1.120 ;
  LAYER metal3 ;
  RECT 1376.800 0.000 1380.340 1.120 ;
  LAYER metal2 ;
  RECT 1376.800 0.000 1380.340 1.120 ;
  LAYER metal1 ;
  RECT 1376.800 0.000 1380.340 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1363.160 0.000 1366.700 1.120 ;
  LAYER metal4 ;
  RECT 1363.160 0.000 1366.700 1.120 ;
  LAYER metal3 ;
  RECT 1363.160 0.000 1366.700 1.120 ;
  LAYER metal2 ;
  RECT 1363.160 0.000 1366.700 1.120 ;
  LAYER metal1 ;
  RECT 1363.160 0.000 1366.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1350.140 0.000 1353.680 1.120 ;
  LAYER metal4 ;
  RECT 1350.140 0.000 1353.680 1.120 ;
  LAYER metal3 ;
  RECT 1350.140 0.000 1353.680 1.120 ;
  LAYER metal2 ;
  RECT 1350.140 0.000 1353.680 1.120 ;
  LAYER metal1 ;
  RECT 1350.140 0.000 1353.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1282.560 0.000 1286.100 1.120 ;
  LAYER metal4 ;
  RECT 1282.560 0.000 1286.100 1.120 ;
  LAYER metal3 ;
  RECT 1282.560 0.000 1286.100 1.120 ;
  LAYER metal2 ;
  RECT 1282.560 0.000 1286.100 1.120 ;
  LAYER metal1 ;
  RECT 1282.560 0.000 1286.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1268.920 0.000 1272.460 1.120 ;
  LAYER metal4 ;
  RECT 1268.920 0.000 1272.460 1.120 ;
  LAYER metal3 ;
  RECT 1268.920 0.000 1272.460 1.120 ;
  LAYER metal2 ;
  RECT 1268.920 0.000 1272.460 1.120 ;
  LAYER metal1 ;
  RECT 1268.920 0.000 1272.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1255.900 0.000 1259.440 1.120 ;
  LAYER metal4 ;
  RECT 1255.900 0.000 1259.440 1.120 ;
  LAYER metal3 ;
  RECT 1255.900 0.000 1259.440 1.120 ;
  LAYER metal2 ;
  RECT 1255.900 0.000 1259.440 1.120 ;
  LAYER metal1 ;
  RECT 1255.900 0.000 1259.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1242.260 0.000 1245.800 1.120 ;
  LAYER metal4 ;
  RECT 1242.260 0.000 1245.800 1.120 ;
  LAYER metal3 ;
  RECT 1242.260 0.000 1245.800 1.120 ;
  LAYER metal2 ;
  RECT 1242.260 0.000 1245.800 1.120 ;
  LAYER metal1 ;
  RECT 1242.260 0.000 1245.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1228.620 0.000 1232.160 1.120 ;
  LAYER metal4 ;
  RECT 1228.620 0.000 1232.160 1.120 ;
  LAYER metal3 ;
  RECT 1228.620 0.000 1232.160 1.120 ;
  LAYER metal2 ;
  RECT 1228.620 0.000 1232.160 1.120 ;
  LAYER metal1 ;
  RECT 1228.620 0.000 1232.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1215.600 0.000 1219.140 1.120 ;
  LAYER metal4 ;
  RECT 1215.600 0.000 1219.140 1.120 ;
  LAYER metal3 ;
  RECT 1215.600 0.000 1219.140 1.120 ;
  LAYER metal2 ;
  RECT 1215.600 0.000 1219.140 1.120 ;
  LAYER metal1 ;
  RECT 1215.600 0.000 1219.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1148.020 0.000 1151.560 1.120 ;
  LAYER metal4 ;
  RECT 1148.020 0.000 1151.560 1.120 ;
  LAYER metal3 ;
  RECT 1148.020 0.000 1151.560 1.120 ;
  LAYER metal2 ;
  RECT 1148.020 0.000 1151.560 1.120 ;
  LAYER metal1 ;
  RECT 1148.020 0.000 1151.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1135.000 0.000 1138.540 1.120 ;
  LAYER metal4 ;
  RECT 1135.000 0.000 1138.540 1.120 ;
  LAYER metal3 ;
  RECT 1135.000 0.000 1138.540 1.120 ;
  LAYER metal2 ;
  RECT 1135.000 0.000 1138.540 1.120 ;
  LAYER metal1 ;
  RECT 1135.000 0.000 1138.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1121.360 0.000 1124.900 1.120 ;
  LAYER metal4 ;
  RECT 1121.360 0.000 1124.900 1.120 ;
  LAYER metal3 ;
  RECT 1121.360 0.000 1124.900 1.120 ;
  LAYER metal2 ;
  RECT 1121.360 0.000 1124.900 1.120 ;
  LAYER metal1 ;
  RECT 1121.360 0.000 1124.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1107.720 0.000 1111.260 1.120 ;
  LAYER metal4 ;
  RECT 1107.720 0.000 1111.260 1.120 ;
  LAYER metal3 ;
  RECT 1107.720 0.000 1111.260 1.120 ;
  LAYER metal2 ;
  RECT 1107.720 0.000 1111.260 1.120 ;
  LAYER metal1 ;
  RECT 1107.720 0.000 1111.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1094.700 0.000 1098.240 1.120 ;
  LAYER metal4 ;
  RECT 1094.700 0.000 1098.240 1.120 ;
  LAYER metal3 ;
  RECT 1094.700 0.000 1098.240 1.120 ;
  LAYER metal2 ;
  RECT 1094.700 0.000 1098.240 1.120 ;
  LAYER metal1 ;
  RECT 1094.700 0.000 1098.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1081.060 0.000 1084.600 1.120 ;
  LAYER metal4 ;
  RECT 1081.060 0.000 1084.600 1.120 ;
  LAYER metal3 ;
  RECT 1081.060 0.000 1084.600 1.120 ;
  LAYER metal2 ;
  RECT 1081.060 0.000 1084.600 1.120 ;
  LAYER metal1 ;
  RECT 1081.060 0.000 1084.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1014.100 0.000 1017.640 1.120 ;
  LAYER metal4 ;
  RECT 1014.100 0.000 1017.640 1.120 ;
  LAYER metal3 ;
  RECT 1014.100 0.000 1017.640 1.120 ;
  LAYER metal2 ;
  RECT 1014.100 0.000 1017.640 1.120 ;
  LAYER metal1 ;
  RECT 1014.100 0.000 1017.640 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1000.460 0.000 1004.000 1.120 ;
  LAYER metal4 ;
  RECT 1000.460 0.000 1004.000 1.120 ;
  LAYER metal3 ;
  RECT 1000.460 0.000 1004.000 1.120 ;
  LAYER metal2 ;
  RECT 1000.460 0.000 1004.000 1.120 ;
  LAYER metal1 ;
  RECT 1000.460 0.000 1004.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 986.820 0.000 990.360 1.120 ;
  LAYER metal4 ;
  RECT 986.820 0.000 990.360 1.120 ;
  LAYER metal3 ;
  RECT 986.820 0.000 990.360 1.120 ;
  LAYER metal2 ;
  RECT 986.820 0.000 990.360 1.120 ;
  LAYER metal1 ;
  RECT 986.820 0.000 990.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 973.800 0.000 977.340 1.120 ;
  LAYER metal4 ;
  RECT 973.800 0.000 977.340 1.120 ;
  LAYER metal3 ;
  RECT 973.800 0.000 977.340 1.120 ;
  LAYER metal2 ;
  RECT 973.800 0.000 977.340 1.120 ;
  LAYER metal1 ;
  RECT 973.800 0.000 977.340 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 960.160 0.000 963.700 1.120 ;
  LAYER metal4 ;
  RECT 960.160 0.000 963.700 1.120 ;
  LAYER metal3 ;
  RECT 960.160 0.000 963.700 1.120 ;
  LAYER metal2 ;
  RECT 960.160 0.000 963.700 1.120 ;
  LAYER metal1 ;
  RECT 960.160 0.000 963.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 946.520 0.000 950.060 1.120 ;
  LAYER metal4 ;
  RECT 946.520 0.000 950.060 1.120 ;
  LAYER metal3 ;
  RECT 946.520 0.000 950.060 1.120 ;
  LAYER metal2 ;
  RECT 946.520 0.000 950.060 1.120 ;
  LAYER metal1 ;
  RECT 946.520 0.000 950.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 881.420 0.000 884.960 1.120 ;
  LAYER metal4 ;
  RECT 881.420 0.000 884.960 1.120 ;
  LAYER metal3 ;
  RECT 881.420 0.000 884.960 1.120 ;
  LAYER metal2 ;
  RECT 881.420 0.000 884.960 1.120 ;
  LAYER metal1 ;
  RECT 881.420 0.000 884.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 865.920 0.000 869.460 1.120 ;
  LAYER metal4 ;
  RECT 865.920 0.000 869.460 1.120 ;
  LAYER metal3 ;
  RECT 865.920 0.000 869.460 1.120 ;
  LAYER metal2 ;
  RECT 865.920 0.000 869.460 1.120 ;
  LAYER metal1 ;
  RECT 865.920 0.000 869.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 852.280 0.000 855.820 1.120 ;
  LAYER metal4 ;
  RECT 852.280 0.000 855.820 1.120 ;
  LAYER metal3 ;
  RECT 852.280 0.000 855.820 1.120 ;
  LAYER metal2 ;
  RECT 852.280 0.000 855.820 1.120 ;
  LAYER metal1 ;
  RECT 852.280 0.000 855.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 839.260 0.000 842.800 1.120 ;
  LAYER metal4 ;
  RECT 839.260 0.000 842.800 1.120 ;
  LAYER metal3 ;
  RECT 839.260 0.000 842.800 1.120 ;
  LAYER metal2 ;
  RECT 839.260 0.000 842.800 1.120 ;
  LAYER metal1 ;
  RECT 839.260 0.000 842.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 825.620 0.000 829.160 1.120 ;
  LAYER metal4 ;
  RECT 825.620 0.000 829.160 1.120 ;
  LAYER metal3 ;
  RECT 825.620 0.000 829.160 1.120 ;
  LAYER metal2 ;
  RECT 825.620 0.000 829.160 1.120 ;
  LAYER metal1 ;
  RECT 825.620 0.000 829.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 811.980 0.000 815.520 1.120 ;
  LAYER metal4 ;
  RECT 811.980 0.000 815.520 1.120 ;
  LAYER metal3 ;
  RECT 811.980 0.000 815.520 1.120 ;
  LAYER metal2 ;
  RECT 811.980 0.000 815.520 1.120 ;
  LAYER metal1 ;
  RECT 811.980 0.000 815.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 745.020 0.000 748.560 1.120 ;
  LAYER metal4 ;
  RECT 745.020 0.000 748.560 1.120 ;
  LAYER metal3 ;
  RECT 745.020 0.000 748.560 1.120 ;
  LAYER metal2 ;
  RECT 745.020 0.000 748.560 1.120 ;
  LAYER metal1 ;
  RECT 745.020 0.000 748.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 731.380 0.000 734.920 1.120 ;
  LAYER metal4 ;
  RECT 731.380 0.000 734.920 1.120 ;
  LAYER metal3 ;
  RECT 731.380 0.000 734.920 1.120 ;
  LAYER metal2 ;
  RECT 731.380 0.000 734.920 1.120 ;
  LAYER metal1 ;
  RECT 731.380 0.000 734.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 718.360 0.000 721.900 1.120 ;
  LAYER metal4 ;
  RECT 718.360 0.000 721.900 1.120 ;
  LAYER metal3 ;
  RECT 718.360 0.000 721.900 1.120 ;
  LAYER metal2 ;
  RECT 718.360 0.000 721.900 1.120 ;
  LAYER metal1 ;
  RECT 718.360 0.000 721.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 704.720 0.000 708.260 1.120 ;
  LAYER metal4 ;
  RECT 704.720 0.000 708.260 1.120 ;
  LAYER metal3 ;
  RECT 704.720 0.000 708.260 1.120 ;
  LAYER metal2 ;
  RECT 704.720 0.000 708.260 1.120 ;
  LAYER metal1 ;
  RECT 704.720 0.000 708.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 691.080 0.000 694.620 1.120 ;
  LAYER metal4 ;
  RECT 691.080 0.000 694.620 1.120 ;
  LAYER metal3 ;
  RECT 691.080 0.000 694.620 1.120 ;
  LAYER metal2 ;
  RECT 691.080 0.000 694.620 1.120 ;
  LAYER metal1 ;
  RECT 691.080 0.000 694.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 678.060 0.000 681.600 1.120 ;
  LAYER metal4 ;
  RECT 678.060 0.000 681.600 1.120 ;
  LAYER metal3 ;
  RECT 678.060 0.000 681.600 1.120 ;
  LAYER metal2 ;
  RECT 678.060 0.000 681.600 1.120 ;
  LAYER metal1 ;
  RECT 678.060 0.000 681.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 610.480 0.000 614.020 1.120 ;
  LAYER metal4 ;
  RECT 610.480 0.000 614.020 1.120 ;
  LAYER metal3 ;
  RECT 610.480 0.000 614.020 1.120 ;
  LAYER metal2 ;
  RECT 610.480 0.000 614.020 1.120 ;
  LAYER metal1 ;
  RECT 610.480 0.000 614.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 597.460 0.000 601.000 1.120 ;
  LAYER metal4 ;
  RECT 597.460 0.000 601.000 1.120 ;
  LAYER metal3 ;
  RECT 597.460 0.000 601.000 1.120 ;
  LAYER metal2 ;
  RECT 597.460 0.000 601.000 1.120 ;
  LAYER metal1 ;
  RECT 597.460 0.000 601.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 583.820 0.000 587.360 1.120 ;
  LAYER metal4 ;
  RECT 583.820 0.000 587.360 1.120 ;
  LAYER metal3 ;
  RECT 583.820 0.000 587.360 1.120 ;
  LAYER metal2 ;
  RECT 583.820 0.000 587.360 1.120 ;
  LAYER metal1 ;
  RECT 583.820 0.000 587.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 570.180 0.000 573.720 1.120 ;
  LAYER metal4 ;
  RECT 570.180 0.000 573.720 1.120 ;
  LAYER metal3 ;
  RECT 570.180 0.000 573.720 1.120 ;
  LAYER metal2 ;
  RECT 570.180 0.000 573.720 1.120 ;
  LAYER metal1 ;
  RECT 570.180 0.000 573.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 557.160 0.000 560.700 1.120 ;
  LAYER metal4 ;
  RECT 557.160 0.000 560.700 1.120 ;
  LAYER metal3 ;
  RECT 557.160 0.000 560.700 1.120 ;
  LAYER metal2 ;
  RECT 557.160 0.000 560.700 1.120 ;
  LAYER metal1 ;
  RECT 557.160 0.000 560.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 543.520 0.000 547.060 1.120 ;
  LAYER metal4 ;
  RECT 543.520 0.000 547.060 1.120 ;
  LAYER metal3 ;
  RECT 543.520 0.000 547.060 1.120 ;
  LAYER metal2 ;
  RECT 543.520 0.000 547.060 1.120 ;
  LAYER metal1 ;
  RECT 543.520 0.000 547.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 475.940 0.000 479.480 1.120 ;
  LAYER metal4 ;
  RECT 475.940 0.000 479.480 1.120 ;
  LAYER metal3 ;
  RECT 475.940 0.000 479.480 1.120 ;
  LAYER metal2 ;
  RECT 475.940 0.000 479.480 1.120 ;
  LAYER metal1 ;
  RECT 475.940 0.000 479.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 462.920 0.000 466.460 1.120 ;
  LAYER metal4 ;
  RECT 462.920 0.000 466.460 1.120 ;
  LAYER metal3 ;
  RECT 462.920 0.000 466.460 1.120 ;
  LAYER metal2 ;
  RECT 462.920 0.000 466.460 1.120 ;
  LAYER metal1 ;
  RECT 462.920 0.000 466.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 451.760 0.000 455.300 1.120 ;
  LAYER metal4 ;
  RECT 451.760 0.000 455.300 1.120 ;
  LAYER metal3 ;
  RECT 451.760 0.000 455.300 1.120 ;
  LAYER metal2 ;
  RECT 451.760 0.000 455.300 1.120 ;
  LAYER metal1 ;
  RECT 451.760 0.000 455.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER metal4 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER metal3 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER metal2 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER metal1 ;
  RECT 435.640 0.000 439.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 422.620 0.000 426.160 1.120 ;
  LAYER metal4 ;
  RECT 422.620 0.000 426.160 1.120 ;
  LAYER metal3 ;
  RECT 422.620 0.000 426.160 1.120 ;
  LAYER metal2 ;
  RECT 422.620 0.000 426.160 1.120 ;
  LAYER metal1 ;
  RECT 422.620 0.000 426.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 408.980 0.000 412.520 1.120 ;
  LAYER metal4 ;
  RECT 408.980 0.000 412.520 1.120 ;
  LAYER metal3 ;
  RECT 408.980 0.000 412.520 1.120 ;
  LAYER metal2 ;
  RECT 408.980 0.000 412.520 1.120 ;
  LAYER metal1 ;
  RECT 408.980 0.000 412.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 342.020 0.000 345.560 1.120 ;
  LAYER metal4 ;
  RECT 342.020 0.000 345.560 1.120 ;
  LAYER metal3 ;
  RECT 342.020 0.000 345.560 1.120 ;
  LAYER metal2 ;
  RECT 342.020 0.000 345.560 1.120 ;
  LAYER metal1 ;
  RECT 342.020 0.000 345.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER metal4 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER metal3 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER metal2 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER metal1 ;
  RECT 328.380 0.000 331.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 314.740 0.000 318.280 1.120 ;
  LAYER metal4 ;
  RECT 314.740 0.000 318.280 1.120 ;
  LAYER metal3 ;
  RECT 314.740 0.000 318.280 1.120 ;
  LAYER metal2 ;
  RECT 314.740 0.000 318.280 1.120 ;
  LAYER metal1 ;
  RECT 314.740 0.000 318.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 301.720 0.000 305.260 1.120 ;
  LAYER metal4 ;
  RECT 301.720 0.000 305.260 1.120 ;
  LAYER metal3 ;
  RECT 301.720 0.000 305.260 1.120 ;
  LAYER metal2 ;
  RECT 301.720 0.000 305.260 1.120 ;
  LAYER metal1 ;
  RECT 301.720 0.000 305.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 288.080 0.000 291.620 1.120 ;
  LAYER metal4 ;
  RECT 288.080 0.000 291.620 1.120 ;
  LAYER metal3 ;
  RECT 288.080 0.000 291.620 1.120 ;
  LAYER metal2 ;
  RECT 288.080 0.000 291.620 1.120 ;
  LAYER metal1 ;
  RECT 288.080 0.000 291.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER metal4 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER metal3 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER metal2 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER metal1 ;
  RECT 274.440 0.000 277.980 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 207.480 0.000 211.020 1.120 ;
  LAYER metal4 ;
  RECT 207.480 0.000 211.020 1.120 ;
  LAYER metal3 ;
  RECT 207.480 0.000 211.020 1.120 ;
  LAYER metal2 ;
  RECT 207.480 0.000 211.020 1.120 ;
  LAYER metal1 ;
  RECT 207.480 0.000 211.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 193.840 0.000 197.380 1.120 ;
  LAYER metal4 ;
  RECT 193.840 0.000 197.380 1.120 ;
  LAYER metal3 ;
  RECT 193.840 0.000 197.380 1.120 ;
  LAYER metal2 ;
  RECT 193.840 0.000 197.380 1.120 ;
  LAYER metal1 ;
  RECT 193.840 0.000 197.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 180.820 0.000 184.360 1.120 ;
  LAYER metal4 ;
  RECT 180.820 0.000 184.360 1.120 ;
  LAYER metal3 ;
  RECT 180.820 0.000 184.360 1.120 ;
  LAYER metal2 ;
  RECT 180.820 0.000 184.360 1.120 ;
  LAYER metal1 ;
  RECT 180.820 0.000 184.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 167.180 0.000 170.720 1.120 ;
  LAYER metal4 ;
  RECT 167.180 0.000 170.720 1.120 ;
  LAYER metal3 ;
  RECT 167.180 0.000 170.720 1.120 ;
  LAYER metal2 ;
  RECT 167.180 0.000 170.720 1.120 ;
  LAYER metal1 ;
  RECT 167.180 0.000 170.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 153.540 0.000 157.080 1.120 ;
  LAYER metal4 ;
  RECT 153.540 0.000 157.080 1.120 ;
  LAYER metal3 ;
  RECT 153.540 0.000 157.080 1.120 ;
  LAYER metal2 ;
  RECT 153.540 0.000 157.080 1.120 ;
  LAYER metal1 ;
  RECT 153.540 0.000 157.080 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER metal4 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER metal3 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER metal2 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER metal1 ;
  RECT 140.520 0.000 144.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 72.940 0.000 76.480 1.120 ;
  LAYER metal4 ;
  RECT 72.940 0.000 76.480 1.120 ;
  LAYER metal3 ;
  RECT 72.940 0.000 76.480 1.120 ;
  LAYER metal2 ;
  RECT 72.940 0.000 76.480 1.120 ;
  LAYER metal1 ;
  RECT 72.940 0.000 76.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER metal4 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER metal3 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER metal2 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER metal1 ;
  RECT 59.300 0.000 62.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER metal4 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER metal3 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER metal2 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER metal1 ;
  RECT 46.280 0.000 49.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER metal4 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER metal3 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER metal2 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER metal1 ;
  RECT 32.640 0.000 36.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 21.480 0.000 25.020 1.120 ;
  LAYER metal4 ;
  RECT 21.480 0.000 25.020 1.120 ;
  LAYER metal3 ;
  RECT 21.480 0.000 25.020 1.120 ;
  LAYER metal2 ;
  RECT 21.480 0.000 25.020 1.120 ;
  LAYER metal1 ;
  RECT 21.480 0.000 25.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER metal4 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER metal3 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER metal2 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER metal1 ;
  RECT 7.220 0.000 10.760 1.120 ;
 END
END VCC
PIN DIB127
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3524.760 178.640 3525.880 179.760 ;
  LAYER metal4 ;
  RECT 3524.760 178.640 3525.880 179.760 ;
  LAYER metal3 ;
  RECT 3524.760 178.640 3525.880 179.760 ;
  LAYER metal2 ;
  RECT 3524.760 178.640 3525.880 179.760 ;
  LAYER metal1 ;
  RECT 3524.760 178.640 3525.880 179.760 ;
 END
END DIB127
PIN DOB127
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3511.120 178.640 3512.240 179.760 ;
  LAYER metal4 ;
  RECT 3511.120 178.640 3512.240 179.760 ;
  LAYER metal3 ;
  RECT 3511.120 178.640 3512.240 179.760 ;
  LAYER metal2 ;
  RECT 3511.120 178.640 3512.240 179.760 ;
  LAYER metal1 ;
  RECT 3511.120 178.640 3512.240 179.760 ;
 END
END DOB127
PIN DIB126
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3497.480 178.640 3498.600 179.760 ;
  LAYER metal4 ;
  RECT 3497.480 178.640 3498.600 179.760 ;
  LAYER metal3 ;
  RECT 3497.480 178.640 3498.600 179.760 ;
  LAYER metal2 ;
  RECT 3497.480 178.640 3498.600 179.760 ;
  LAYER metal1 ;
  RECT 3497.480 178.640 3498.600 179.760 ;
 END
END DIB126
PIN DOB126
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3484.460 178.640 3485.580 179.760 ;
  LAYER metal4 ;
  RECT 3484.460 178.640 3485.580 179.760 ;
  LAYER metal3 ;
  RECT 3484.460 178.640 3485.580 179.760 ;
  LAYER metal2 ;
  RECT 3484.460 178.640 3485.580 179.760 ;
  LAYER metal1 ;
  RECT 3484.460 178.640 3485.580 179.760 ;
 END
END DOB126
PIN DIB125
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3470.820 178.640 3471.940 179.760 ;
  LAYER metal4 ;
  RECT 3470.820 178.640 3471.940 179.760 ;
  LAYER metal3 ;
  RECT 3470.820 178.640 3471.940 179.760 ;
  LAYER metal2 ;
  RECT 3470.820 178.640 3471.940 179.760 ;
  LAYER metal1 ;
  RECT 3470.820 178.640 3471.940 179.760 ;
 END
END DIB125
PIN DOB125
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3457.180 178.640 3458.300 179.760 ;
  LAYER metal4 ;
  RECT 3457.180 178.640 3458.300 179.760 ;
  LAYER metal3 ;
  RECT 3457.180 178.640 3458.300 179.760 ;
  LAYER metal2 ;
  RECT 3457.180 178.640 3458.300 179.760 ;
  LAYER metal1 ;
  RECT 3457.180 178.640 3458.300 179.760 ;
 END
END DOB125
PIN DIB124
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3444.160 178.640 3445.280 179.760 ;
  LAYER metal4 ;
  RECT 3444.160 178.640 3445.280 179.760 ;
  LAYER metal3 ;
  RECT 3444.160 178.640 3445.280 179.760 ;
  LAYER metal2 ;
  RECT 3444.160 178.640 3445.280 179.760 ;
  LAYER metal1 ;
  RECT 3444.160 178.640 3445.280 179.760 ;
 END
END DIB124
PIN DOB124
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3430.520 178.640 3431.640 179.760 ;
  LAYER metal4 ;
  RECT 3430.520 178.640 3431.640 179.760 ;
  LAYER metal3 ;
  RECT 3430.520 178.640 3431.640 179.760 ;
  LAYER metal2 ;
  RECT 3430.520 178.640 3431.640 179.760 ;
  LAYER metal1 ;
  RECT 3430.520 178.640 3431.640 179.760 ;
 END
END DOB124
PIN DIB123
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3416.880 178.640 3418.000 179.760 ;
  LAYER metal4 ;
  RECT 3416.880 178.640 3418.000 179.760 ;
  LAYER metal3 ;
  RECT 3416.880 178.640 3418.000 179.760 ;
  LAYER metal2 ;
  RECT 3416.880 178.640 3418.000 179.760 ;
  LAYER metal1 ;
  RECT 3416.880 178.640 3418.000 179.760 ;
 END
END DIB123
PIN DOB123
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3403.860 178.640 3404.980 179.760 ;
  LAYER metal4 ;
  RECT 3403.860 178.640 3404.980 179.760 ;
  LAYER metal3 ;
  RECT 3403.860 178.640 3404.980 179.760 ;
  LAYER metal2 ;
  RECT 3403.860 178.640 3404.980 179.760 ;
  LAYER metal1 ;
  RECT 3403.860 178.640 3404.980 179.760 ;
 END
END DOB123
PIN DIB122
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3390.220 178.640 3391.340 179.760 ;
  LAYER metal4 ;
  RECT 3390.220 178.640 3391.340 179.760 ;
  LAYER metal3 ;
  RECT 3390.220 178.640 3391.340 179.760 ;
  LAYER metal2 ;
  RECT 3390.220 178.640 3391.340 179.760 ;
  LAYER metal1 ;
  RECT 3390.220 178.640 3391.340 179.760 ;
 END
END DIB122
PIN DOB122
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3376.580 178.640 3377.700 179.760 ;
  LAYER metal4 ;
  RECT 3376.580 178.640 3377.700 179.760 ;
  LAYER metal3 ;
  RECT 3376.580 178.640 3377.700 179.760 ;
  LAYER metal2 ;
  RECT 3376.580 178.640 3377.700 179.760 ;
  LAYER metal1 ;
  RECT 3376.580 178.640 3377.700 179.760 ;
 END
END DOB122
PIN DIB121
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3363.560 178.640 3364.680 179.760 ;
  LAYER metal4 ;
  RECT 3363.560 178.640 3364.680 179.760 ;
  LAYER metal3 ;
  RECT 3363.560 178.640 3364.680 179.760 ;
  LAYER metal2 ;
  RECT 3363.560 178.640 3364.680 179.760 ;
  LAYER metal1 ;
  RECT 3363.560 178.640 3364.680 179.760 ;
 END
END DIB121
PIN DOB121
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3349.920 178.640 3351.040 179.760 ;
  LAYER metal4 ;
  RECT 3349.920 178.640 3351.040 179.760 ;
  LAYER metal3 ;
  RECT 3349.920 178.640 3351.040 179.760 ;
  LAYER metal2 ;
  RECT 3349.920 178.640 3351.040 179.760 ;
  LAYER metal1 ;
  RECT 3349.920 178.640 3351.040 179.760 ;
 END
END DOB121
PIN DIB120
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3336.280 178.640 3337.400 179.760 ;
  LAYER metal4 ;
  RECT 3336.280 178.640 3337.400 179.760 ;
  LAYER metal3 ;
  RECT 3336.280 178.640 3337.400 179.760 ;
  LAYER metal2 ;
  RECT 3336.280 178.640 3337.400 179.760 ;
  LAYER metal1 ;
  RECT 3336.280 178.640 3337.400 179.760 ;
 END
END DIB120
PIN DOB120
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3322.640 178.640 3323.760 179.760 ;
  LAYER metal4 ;
  RECT 3322.640 178.640 3323.760 179.760 ;
  LAYER metal3 ;
  RECT 3322.640 178.640 3323.760 179.760 ;
  LAYER metal2 ;
  RECT 3322.640 178.640 3323.760 179.760 ;
  LAYER metal1 ;
  RECT 3322.640 178.640 3323.760 179.760 ;
 END
END DOB120
PIN DIB119
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3309.620 178.640 3310.740 179.760 ;
  LAYER metal4 ;
  RECT 3309.620 178.640 3310.740 179.760 ;
  LAYER metal3 ;
  RECT 3309.620 178.640 3310.740 179.760 ;
  LAYER metal2 ;
  RECT 3309.620 178.640 3310.740 179.760 ;
  LAYER metal1 ;
  RECT 3309.620 178.640 3310.740 179.760 ;
 END
END DIB119
PIN DOB119
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3295.980 178.640 3297.100 179.760 ;
  LAYER metal4 ;
  RECT 3295.980 178.640 3297.100 179.760 ;
  LAYER metal3 ;
  RECT 3295.980 178.640 3297.100 179.760 ;
  LAYER metal2 ;
  RECT 3295.980 178.640 3297.100 179.760 ;
  LAYER metal1 ;
  RECT 3295.980 178.640 3297.100 179.760 ;
 END
END DOB119
PIN DIB118
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3282.340 178.640 3283.460 179.760 ;
  LAYER metal4 ;
  RECT 3282.340 178.640 3283.460 179.760 ;
  LAYER metal3 ;
  RECT 3282.340 178.640 3283.460 179.760 ;
  LAYER metal2 ;
  RECT 3282.340 178.640 3283.460 179.760 ;
  LAYER metal1 ;
  RECT 3282.340 178.640 3283.460 179.760 ;
 END
END DIB118
PIN DOB118
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3269.320 178.640 3270.440 179.760 ;
  LAYER metal4 ;
  RECT 3269.320 178.640 3270.440 179.760 ;
  LAYER metal3 ;
  RECT 3269.320 178.640 3270.440 179.760 ;
  LAYER metal2 ;
  RECT 3269.320 178.640 3270.440 179.760 ;
  LAYER metal1 ;
  RECT 3269.320 178.640 3270.440 179.760 ;
 END
END DOB118
PIN DIB117
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3255.680 178.640 3256.800 179.760 ;
  LAYER metal4 ;
  RECT 3255.680 178.640 3256.800 179.760 ;
  LAYER metal3 ;
  RECT 3255.680 178.640 3256.800 179.760 ;
  LAYER metal2 ;
  RECT 3255.680 178.640 3256.800 179.760 ;
  LAYER metal1 ;
  RECT 3255.680 178.640 3256.800 179.760 ;
 END
END DIB117
PIN DOB117
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3242.040 178.640 3243.160 179.760 ;
  LAYER metal4 ;
  RECT 3242.040 178.640 3243.160 179.760 ;
  LAYER metal3 ;
  RECT 3242.040 178.640 3243.160 179.760 ;
  LAYER metal2 ;
  RECT 3242.040 178.640 3243.160 179.760 ;
  LAYER metal1 ;
  RECT 3242.040 178.640 3243.160 179.760 ;
 END
END DOB117
PIN DIB116
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3229.020 178.640 3230.140 179.760 ;
  LAYER metal4 ;
  RECT 3229.020 178.640 3230.140 179.760 ;
  LAYER metal3 ;
  RECT 3229.020 178.640 3230.140 179.760 ;
  LAYER metal2 ;
  RECT 3229.020 178.640 3230.140 179.760 ;
  LAYER metal1 ;
  RECT 3229.020 178.640 3230.140 179.760 ;
 END
END DIB116
PIN DOB116
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3215.380 178.640 3216.500 179.760 ;
  LAYER metal4 ;
  RECT 3215.380 178.640 3216.500 179.760 ;
  LAYER metal3 ;
  RECT 3215.380 178.640 3216.500 179.760 ;
  LAYER metal2 ;
  RECT 3215.380 178.640 3216.500 179.760 ;
  LAYER metal1 ;
  RECT 3215.380 178.640 3216.500 179.760 ;
 END
END DOB116
PIN DIB115
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3201.740 178.640 3202.860 179.760 ;
  LAYER metal4 ;
  RECT 3201.740 178.640 3202.860 179.760 ;
  LAYER metal3 ;
  RECT 3201.740 178.640 3202.860 179.760 ;
  LAYER metal2 ;
  RECT 3201.740 178.640 3202.860 179.760 ;
  LAYER metal1 ;
  RECT 3201.740 178.640 3202.860 179.760 ;
 END
END DIB115
PIN DOB115
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3188.720 178.640 3189.840 179.760 ;
  LAYER metal4 ;
  RECT 3188.720 178.640 3189.840 179.760 ;
  LAYER metal3 ;
  RECT 3188.720 178.640 3189.840 179.760 ;
  LAYER metal2 ;
  RECT 3188.720 178.640 3189.840 179.760 ;
  LAYER metal1 ;
  RECT 3188.720 178.640 3189.840 179.760 ;
 END
END DOB115
PIN DIB114
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3175.080 178.640 3176.200 179.760 ;
  LAYER metal4 ;
  RECT 3175.080 178.640 3176.200 179.760 ;
  LAYER metal3 ;
  RECT 3175.080 178.640 3176.200 179.760 ;
  LAYER metal2 ;
  RECT 3175.080 178.640 3176.200 179.760 ;
  LAYER metal1 ;
  RECT 3175.080 178.640 3176.200 179.760 ;
 END
END DIB114
PIN DOB114
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3161.440 178.640 3162.560 179.760 ;
  LAYER metal4 ;
  RECT 3161.440 178.640 3162.560 179.760 ;
  LAYER metal3 ;
  RECT 3161.440 178.640 3162.560 179.760 ;
  LAYER metal2 ;
  RECT 3161.440 178.640 3162.560 179.760 ;
  LAYER metal1 ;
  RECT 3161.440 178.640 3162.560 179.760 ;
 END
END DOB114
PIN DIB113
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3148.420 178.640 3149.540 179.760 ;
  LAYER metal4 ;
  RECT 3148.420 178.640 3149.540 179.760 ;
  LAYER metal3 ;
  RECT 3148.420 178.640 3149.540 179.760 ;
  LAYER metal2 ;
  RECT 3148.420 178.640 3149.540 179.760 ;
  LAYER metal1 ;
  RECT 3148.420 178.640 3149.540 179.760 ;
 END
END DIB113
PIN DOB113
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3134.780 178.640 3135.900 179.760 ;
  LAYER metal4 ;
  RECT 3134.780 178.640 3135.900 179.760 ;
  LAYER metal3 ;
  RECT 3134.780 178.640 3135.900 179.760 ;
  LAYER metal2 ;
  RECT 3134.780 178.640 3135.900 179.760 ;
  LAYER metal1 ;
  RECT 3134.780 178.640 3135.900 179.760 ;
 END
END DOB113
PIN DIB112
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3121.140 178.640 3122.260 179.760 ;
  LAYER metal4 ;
  RECT 3121.140 178.640 3122.260 179.760 ;
  LAYER metal3 ;
  RECT 3121.140 178.640 3122.260 179.760 ;
  LAYER metal2 ;
  RECT 3121.140 178.640 3122.260 179.760 ;
  LAYER metal1 ;
  RECT 3121.140 178.640 3122.260 179.760 ;
 END
END DIB112
PIN WEBN7
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3109.980 178.640 3111.100 179.760 ;
  LAYER metal4 ;
  RECT 3109.980 178.640 3111.100 179.760 ;
  LAYER metal3 ;
  RECT 3109.980 178.640 3111.100 179.760 ;
  LAYER metal2 ;
  RECT 3109.980 178.640 3111.100 179.760 ;
  LAYER metal1 ;
  RECT 3109.980 178.640 3111.100 179.760 ;
 END
END WEBN7
PIN DOB112
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3108.120 178.640 3109.240 179.760 ;
  LAYER metal4 ;
  RECT 3108.120 178.640 3109.240 179.760 ;
  LAYER metal3 ;
  RECT 3108.120 178.640 3109.240 179.760 ;
  LAYER metal2 ;
  RECT 3108.120 178.640 3109.240 179.760 ;
  LAYER metal1 ;
  RECT 3108.120 178.640 3109.240 179.760 ;
 END
END DOB112
PIN DIB111
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3094.480 178.640 3095.600 179.760 ;
  LAYER metal4 ;
  RECT 3094.480 178.640 3095.600 179.760 ;
  LAYER metal3 ;
  RECT 3094.480 178.640 3095.600 179.760 ;
  LAYER metal2 ;
  RECT 3094.480 178.640 3095.600 179.760 ;
  LAYER metal1 ;
  RECT 3094.480 178.640 3095.600 179.760 ;
 END
END DIB111
PIN DOB111
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3080.840 178.640 3081.960 179.760 ;
  LAYER metal4 ;
  RECT 3080.840 178.640 3081.960 179.760 ;
  LAYER metal3 ;
  RECT 3080.840 178.640 3081.960 179.760 ;
  LAYER metal2 ;
  RECT 3080.840 178.640 3081.960 179.760 ;
  LAYER metal1 ;
  RECT 3080.840 178.640 3081.960 179.760 ;
 END
END DOB111
PIN DIB110
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3067.820 178.640 3068.940 179.760 ;
  LAYER metal4 ;
  RECT 3067.820 178.640 3068.940 179.760 ;
  LAYER metal3 ;
  RECT 3067.820 178.640 3068.940 179.760 ;
  LAYER metal2 ;
  RECT 3067.820 178.640 3068.940 179.760 ;
  LAYER metal1 ;
  RECT 3067.820 178.640 3068.940 179.760 ;
 END
END DIB110
PIN DOB110
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3054.180 178.640 3055.300 179.760 ;
  LAYER metal4 ;
  RECT 3054.180 178.640 3055.300 179.760 ;
  LAYER metal3 ;
  RECT 3054.180 178.640 3055.300 179.760 ;
  LAYER metal2 ;
  RECT 3054.180 178.640 3055.300 179.760 ;
  LAYER metal1 ;
  RECT 3054.180 178.640 3055.300 179.760 ;
 END
END DOB110
PIN DIB109
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3040.540 178.640 3041.660 179.760 ;
  LAYER metal4 ;
  RECT 3040.540 178.640 3041.660 179.760 ;
  LAYER metal3 ;
  RECT 3040.540 178.640 3041.660 179.760 ;
  LAYER metal2 ;
  RECT 3040.540 178.640 3041.660 179.760 ;
  LAYER metal1 ;
  RECT 3040.540 178.640 3041.660 179.760 ;
 END
END DIB109
PIN DOB109
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3027.520 178.640 3028.640 179.760 ;
  LAYER metal4 ;
  RECT 3027.520 178.640 3028.640 179.760 ;
  LAYER metal3 ;
  RECT 3027.520 178.640 3028.640 179.760 ;
  LAYER metal2 ;
  RECT 3027.520 178.640 3028.640 179.760 ;
  LAYER metal1 ;
  RECT 3027.520 178.640 3028.640 179.760 ;
 END
END DOB109
PIN DIB108
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3013.880 178.640 3015.000 179.760 ;
  LAYER metal4 ;
  RECT 3013.880 178.640 3015.000 179.760 ;
  LAYER metal3 ;
  RECT 3013.880 178.640 3015.000 179.760 ;
  LAYER metal2 ;
  RECT 3013.880 178.640 3015.000 179.760 ;
  LAYER metal1 ;
  RECT 3013.880 178.640 3015.000 179.760 ;
 END
END DIB108
PIN DOB108
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3000.240 178.640 3001.360 179.760 ;
  LAYER metal4 ;
  RECT 3000.240 178.640 3001.360 179.760 ;
  LAYER metal3 ;
  RECT 3000.240 178.640 3001.360 179.760 ;
  LAYER metal2 ;
  RECT 3000.240 178.640 3001.360 179.760 ;
  LAYER metal1 ;
  RECT 3000.240 178.640 3001.360 179.760 ;
 END
END DOB108
PIN DIB107
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2987.220 178.640 2988.340 179.760 ;
  LAYER metal4 ;
  RECT 2987.220 178.640 2988.340 179.760 ;
  LAYER metal3 ;
  RECT 2987.220 178.640 2988.340 179.760 ;
  LAYER metal2 ;
  RECT 2987.220 178.640 2988.340 179.760 ;
  LAYER metal1 ;
  RECT 2987.220 178.640 2988.340 179.760 ;
 END
END DIB107
PIN DOB107
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2973.580 178.640 2974.700 179.760 ;
  LAYER metal4 ;
  RECT 2973.580 178.640 2974.700 179.760 ;
  LAYER metal3 ;
  RECT 2973.580 178.640 2974.700 179.760 ;
  LAYER metal2 ;
  RECT 2973.580 178.640 2974.700 179.760 ;
  LAYER metal1 ;
  RECT 2973.580 178.640 2974.700 179.760 ;
 END
END DOB107
PIN DIB106
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2959.940 178.640 2961.060 179.760 ;
  LAYER metal4 ;
  RECT 2959.940 178.640 2961.060 179.760 ;
  LAYER metal3 ;
  RECT 2959.940 178.640 2961.060 179.760 ;
  LAYER metal2 ;
  RECT 2959.940 178.640 2961.060 179.760 ;
  LAYER metal1 ;
  RECT 2959.940 178.640 2961.060 179.760 ;
 END
END DIB106
PIN DOB106
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2946.920 178.640 2948.040 179.760 ;
  LAYER metal4 ;
  RECT 2946.920 178.640 2948.040 179.760 ;
  LAYER metal3 ;
  RECT 2946.920 178.640 2948.040 179.760 ;
  LAYER metal2 ;
  RECT 2946.920 178.640 2948.040 179.760 ;
  LAYER metal1 ;
  RECT 2946.920 178.640 2948.040 179.760 ;
 END
END DOB106
PIN DIB105
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2933.280 178.640 2934.400 179.760 ;
  LAYER metal4 ;
  RECT 2933.280 178.640 2934.400 179.760 ;
  LAYER metal3 ;
  RECT 2933.280 178.640 2934.400 179.760 ;
  LAYER metal2 ;
  RECT 2933.280 178.640 2934.400 179.760 ;
  LAYER metal1 ;
  RECT 2933.280 178.640 2934.400 179.760 ;
 END
END DIB105
PIN DOB105
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2919.640 178.640 2920.760 179.760 ;
  LAYER metal4 ;
  RECT 2919.640 178.640 2920.760 179.760 ;
  LAYER metal3 ;
  RECT 2919.640 178.640 2920.760 179.760 ;
  LAYER metal2 ;
  RECT 2919.640 178.640 2920.760 179.760 ;
  LAYER metal1 ;
  RECT 2919.640 178.640 2920.760 179.760 ;
 END
END DOB105
PIN DIB104
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2906.000 178.640 2907.120 179.760 ;
  LAYER metal4 ;
  RECT 2906.000 178.640 2907.120 179.760 ;
  LAYER metal3 ;
  RECT 2906.000 178.640 2907.120 179.760 ;
  LAYER metal2 ;
  RECT 2906.000 178.640 2907.120 179.760 ;
  LAYER metal1 ;
  RECT 2906.000 178.640 2907.120 179.760 ;
 END
END DIB104
PIN DOB104
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2892.980 178.640 2894.100 179.760 ;
  LAYER metal4 ;
  RECT 2892.980 178.640 2894.100 179.760 ;
  LAYER metal3 ;
  RECT 2892.980 178.640 2894.100 179.760 ;
  LAYER metal2 ;
  RECT 2892.980 178.640 2894.100 179.760 ;
  LAYER metal1 ;
  RECT 2892.980 178.640 2894.100 179.760 ;
 END
END DOB104
PIN DIB103
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2879.340 178.640 2880.460 179.760 ;
  LAYER metal4 ;
  RECT 2879.340 178.640 2880.460 179.760 ;
  LAYER metal3 ;
  RECT 2879.340 178.640 2880.460 179.760 ;
  LAYER metal2 ;
  RECT 2879.340 178.640 2880.460 179.760 ;
  LAYER metal1 ;
  RECT 2879.340 178.640 2880.460 179.760 ;
 END
END DIB103
PIN DOB103
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2865.700 178.640 2866.820 179.760 ;
  LAYER metal4 ;
  RECT 2865.700 178.640 2866.820 179.760 ;
  LAYER metal3 ;
  RECT 2865.700 178.640 2866.820 179.760 ;
  LAYER metal2 ;
  RECT 2865.700 178.640 2866.820 179.760 ;
  LAYER metal1 ;
  RECT 2865.700 178.640 2866.820 179.760 ;
 END
END DOB103
PIN DIB102
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2852.680 178.640 2853.800 179.760 ;
  LAYER metal4 ;
  RECT 2852.680 178.640 2853.800 179.760 ;
  LAYER metal3 ;
  RECT 2852.680 178.640 2853.800 179.760 ;
  LAYER metal2 ;
  RECT 2852.680 178.640 2853.800 179.760 ;
  LAYER metal1 ;
  RECT 2852.680 178.640 2853.800 179.760 ;
 END
END DIB102
PIN DOB102
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2839.040 178.640 2840.160 179.760 ;
  LAYER metal4 ;
  RECT 2839.040 178.640 2840.160 179.760 ;
  LAYER metal3 ;
  RECT 2839.040 178.640 2840.160 179.760 ;
  LAYER metal2 ;
  RECT 2839.040 178.640 2840.160 179.760 ;
  LAYER metal1 ;
  RECT 2839.040 178.640 2840.160 179.760 ;
 END
END DOB102
PIN DIB101
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2825.400 178.640 2826.520 179.760 ;
  LAYER metal4 ;
  RECT 2825.400 178.640 2826.520 179.760 ;
  LAYER metal3 ;
  RECT 2825.400 178.640 2826.520 179.760 ;
  LAYER metal2 ;
  RECT 2825.400 178.640 2826.520 179.760 ;
  LAYER metal1 ;
  RECT 2825.400 178.640 2826.520 179.760 ;
 END
END DIB101
PIN DOB101
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2812.380 178.640 2813.500 179.760 ;
  LAYER metal4 ;
  RECT 2812.380 178.640 2813.500 179.760 ;
  LAYER metal3 ;
  RECT 2812.380 178.640 2813.500 179.760 ;
  LAYER metal2 ;
  RECT 2812.380 178.640 2813.500 179.760 ;
  LAYER metal1 ;
  RECT 2812.380 178.640 2813.500 179.760 ;
 END
END DOB101
PIN DIB100
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2798.740 178.640 2799.860 179.760 ;
  LAYER metal4 ;
  RECT 2798.740 178.640 2799.860 179.760 ;
  LAYER metal3 ;
  RECT 2798.740 178.640 2799.860 179.760 ;
  LAYER metal2 ;
  RECT 2798.740 178.640 2799.860 179.760 ;
  LAYER metal1 ;
  RECT 2798.740 178.640 2799.860 179.760 ;
 END
END DIB100
PIN DOB100
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2785.100 178.640 2786.220 179.760 ;
  LAYER metal4 ;
  RECT 2785.100 178.640 2786.220 179.760 ;
  LAYER metal3 ;
  RECT 2785.100 178.640 2786.220 179.760 ;
  LAYER metal2 ;
  RECT 2785.100 178.640 2786.220 179.760 ;
  LAYER metal1 ;
  RECT 2785.100 178.640 2786.220 179.760 ;
 END
END DOB100
PIN DIB99
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2772.080 178.640 2773.200 179.760 ;
  LAYER metal4 ;
  RECT 2772.080 178.640 2773.200 179.760 ;
  LAYER metal3 ;
  RECT 2772.080 178.640 2773.200 179.760 ;
  LAYER metal2 ;
  RECT 2772.080 178.640 2773.200 179.760 ;
  LAYER metal1 ;
  RECT 2772.080 178.640 2773.200 179.760 ;
 END
END DIB99
PIN DOB99
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2758.440 178.640 2759.560 179.760 ;
  LAYER metal4 ;
  RECT 2758.440 178.640 2759.560 179.760 ;
  LAYER metal3 ;
  RECT 2758.440 178.640 2759.560 179.760 ;
  LAYER metal2 ;
  RECT 2758.440 178.640 2759.560 179.760 ;
  LAYER metal1 ;
  RECT 2758.440 178.640 2759.560 179.760 ;
 END
END DOB99
PIN DIB98
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2744.800 178.640 2745.920 179.760 ;
  LAYER metal4 ;
  RECT 2744.800 178.640 2745.920 179.760 ;
  LAYER metal3 ;
  RECT 2744.800 178.640 2745.920 179.760 ;
  LAYER metal2 ;
  RECT 2744.800 178.640 2745.920 179.760 ;
  LAYER metal1 ;
  RECT 2744.800 178.640 2745.920 179.760 ;
 END
END DIB98
PIN DOB98
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2731.780 178.640 2732.900 179.760 ;
  LAYER metal4 ;
  RECT 2731.780 178.640 2732.900 179.760 ;
  LAYER metal3 ;
  RECT 2731.780 178.640 2732.900 179.760 ;
  LAYER metal2 ;
  RECT 2731.780 178.640 2732.900 179.760 ;
  LAYER metal1 ;
  RECT 2731.780 178.640 2732.900 179.760 ;
 END
END DOB98
PIN DIB97
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2718.140 178.640 2719.260 179.760 ;
  LAYER metal4 ;
  RECT 2718.140 178.640 2719.260 179.760 ;
  LAYER metal3 ;
  RECT 2718.140 178.640 2719.260 179.760 ;
  LAYER metal2 ;
  RECT 2718.140 178.640 2719.260 179.760 ;
  LAYER metal1 ;
  RECT 2718.140 178.640 2719.260 179.760 ;
 END
END DIB97
PIN DOB97
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2704.500 178.640 2705.620 179.760 ;
  LAYER metal4 ;
  RECT 2704.500 178.640 2705.620 179.760 ;
  LAYER metal3 ;
  RECT 2704.500 178.640 2705.620 179.760 ;
  LAYER metal2 ;
  RECT 2704.500 178.640 2705.620 179.760 ;
  LAYER metal1 ;
  RECT 2704.500 178.640 2705.620 179.760 ;
 END
END DOB97
PIN DIB96
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2691.480 178.640 2692.600 179.760 ;
  LAYER metal4 ;
  RECT 2691.480 178.640 2692.600 179.760 ;
  LAYER metal3 ;
  RECT 2691.480 178.640 2692.600 179.760 ;
  LAYER metal2 ;
  RECT 2691.480 178.640 2692.600 179.760 ;
  LAYER metal1 ;
  RECT 2691.480 178.640 2692.600 179.760 ;
 END
END DIB96
PIN WEBN6
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2680.320 178.640 2681.440 179.760 ;
  LAYER metal4 ;
  RECT 2680.320 178.640 2681.440 179.760 ;
  LAYER metal3 ;
  RECT 2680.320 178.640 2681.440 179.760 ;
  LAYER metal2 ;
  RECT 2680.320 178.640 2681.440 179.760 ;
  LAYER metal1 ;
  RECT 2680.320 178.640 2681.440 179.760 ;
 END
END WEBN6
PIN DOB96
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2677.840 178.640 2678.960 179.760 ;
  LAYER metal4 ;
  RECT 2677.840 178.640 2678.960 179.760 ;
  LAYER metal3 ;
  RECT 2677.840 178.640 2678.960 179.760 ;
  LAYER metal2 ;
  RECT 2677.840 178.640 2678.960 179.760 ;
  LAYER metal1 ;
  RECT 2677.840 178.640 2678.960 179.760 ;
 END
END DOB96
PIN DIB95
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2664.200 178.640 2665.320 179.760 ;
  LAYER metal4 ;
  RECT 2664.200 178.640 2665.320 179.760 ;
  LAYER metal3 ;
  RECT 2664.200 178.640 2665.320 179.760 ;
  LAYER metal2 ;
  RECT 2664.200 178.640 2665.320 179.760 ;
  LAYER metal1 ;
  RECT 2664.200 178.640 2665.320 179.760 ;
 END
END DIB95
PIN DOB95
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2651.180 178.640 2652.300 179.760 ;
  LAYER metal4 ;
  RECT 2651.180 178.640 2652.300 179.760 ;
  LAYER metal3 ;
  RECT 2651.180 178.640 2652.300 179.760 ;
  LAYER metal2 ;
  RECT 2651.180 178.640 2652.300 179.760 ;
  LAYER metal1 ;
  RECT 2651.180 178.640 2652.300 179.760 ;
 END
END DOB95
PIN DIB94
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2637.540 178.640 2638.660 179.760 ;
  LAYER metal4 ;
  RECT 2637.540 178.640 2638.660 179.760 ;
  LAYER metal3 ;
  RECT 2637.540 178.640 2638.660 179.760 ;
  LAYER metal2 ;
  RECT 2637.540 178.640 2638.660 179.760 ;
  LAYER metal1 ;
  RECT 2637.540 178.640 2638.660 179.760 ;
 END
END DIB94
PIN DOB94
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2623.900 178.640 2625.020 179.760 ;
  LAYER metal4 ;
  RECT 2623.900 178.640 2625.020 179.760 ;
  LAYER metal3 ;
  RECT 2623.900 178.640 2625.020 179.760 ;
  LAYER metal2 ;
  RECT 2623.900 178.640 2625.020 179.760 ;
  LAYER metal1 ;
  RECT 2623.900 178.640 2625.020 179.760 ;
 END
END DOB94
PIN DIB93
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2610.880 178.640 2612.000 179.760 ;
  LAYER metal4 ;
  RECT 2610.880 178.640 2612.000 179.760 ;
  LAYER metal3 ;
  RECT 2610.880 178.640 2612.000 179.760 ;
  LAYER metal2 ;
  RECT 2610.880 178.640 2612.000 179.760 ;
  LAYER metal1 ;
  RECT 2610.880 178.640 2612.000 179.760 ;
 END
END DIB93
PIN DOB93
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2597.240 178.640 2598.360 179.760 ;
  LAYER metal4 ;
  RECT 2597.240 178.640 2598.360 179.760 ;
  LAYER metal3 ;
  RECT 2597.240 178.640 2598.360 179.760 ;
  LAYER metal2 ;
  RECT 2597.240 178.640 2598.360 179.760 ;
  LAYER metal1 ;
  RECT 2597.240 178.640 2598.360 179.760 ;
 END
END DOB93
PIN DIB92
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2583.600 178.640 2584.720 179.760 ;
  LAYER metal4 ;
  RECT 2583.600 178.640 2584.720 179.760 ;
  LAYER metal3 ;
  RECT 2583.600 178.640 2584.720 179.760 ;
  LAYER metal2 ;
  RECT 2583.600 178.640 2584.720 179.760 ;
  LAYER metal1 ;
  RECT 2583.600 178.640 2584.720 179.760 ;
 END
END DIB92
PIN DOB92
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2570.580 178.640 2571.700 179.760 ;
  LAYER metal4 ;
  RECT 2570.580 178.640 2571.700 179.760 ;
  LAYER metal3 ;
  RECT 2570.580 178.640 2571.700 179.760 ;
  LAYER metal2 ;
  RECT 2570.580 178.640 2571.700 179.760 ;
  LAYER metal1 ;
  RECT 2570.580 178.640 2571.700 179.760 ;
 END
END DOB92
PIN DIB91
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2556.940 178.640 2558.060 179.760 ;
  LAYER metal4 ;
  RECT 2556.940 178.640 2558.060 179.760 ;
  LAYER metal3 ;
  RECT 2556.940 178.640 2558.060 179.760 ;
  LAYER metal2 ;
  RECT 2556.940 178.640 2558.060 179.760 ;
  LAYER metal1 ;
  RECT 2556.940 178.640 2558.060 179.760 ;
 END
END DIB91
PIN DOB91
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2543.300 178.640 2544.420 179.760 ;
  LAYER metal4 ;
  RECT 2543.300 178.640 2544.420 179.760 ;
  LAYER metal3 ;
  RECT 2543.300 178.640 2544.420 179.760 ;
  LAYER metal2 ;
  RECT 2543.300 178.640 2544.420 179.760 ;
  LAYER metal1 ;
  RECT 2543.300 178.640 2544.420 179.760 ;
 END
END DOB91
PIN DIB90
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2530.280 178.640 2531.400 179.760 ;
  LAYER metal4 ;
  RECT 2530.280 178.640 2531.400 179.760 ;
  LAYER metal3 ;
  RECT 2530.280 178.640 2531.400 179.760 ;
  LAYER metal2 ;
  RECT 2530.280 178.640 2531.400 179.760 ;
  LAYER metal1 ;
  RECT 2530.280 178.640 2531.400 179.760 ;
 END
END DIB90
PIN DOB90
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2516.640 178.640 2517.760 179.760 ;
  LAYER metal4 ;
  RECT 2516.640 178.640 2517.760 179.760 ;
  LAYER metal3 ;
  RECT 2516.640 178.640 2517.760 179.760 ;
  LAYER metal2 ;
  RECT 2516.640 178.640 2517.760 179.760 ;
  LAYER metal1 ;
  RECT 2516.640 178.640 2517.760 179.760 ;
 END
END DOB90
PIN DIB89
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2503.000 178.640 2504.120 179.760 ;
  LAYER metal4 ;
  RECT 2503.000 178.640 2504.120 179.760 ;
  LAYER metal3 ;
  RECT 2503.000 178.640 2504.120 179.760 ;
  LAYER metal2 ;
  RECT 2503.000 178.640 2504.120 179.760 ;
  LAYER metal1 ;
  RECT 2503.000 178.640 2504.120 179.760 ;
 END
END DIB89
PIN DOB89
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2489.360 178.640 2490.480 179.760 ;
  LAYER metal4 ;
  RECT 2489.360 178.640 2490.480 179.760 ;
  LAYER metal3 ;
  RECT 2489.360 178.640 2490.480 179.760 ;
  LAYER metal2 ;
  RECT 2489.360 178.640 2490.480 179.760 ;
  LAYER metal1 ;
  RECT 2489.360 178.640 2490.480 179.760 ;
 END
END DOB89
PIN DIB88
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2476.340 178.640 2477.460 179.760 ;
  LAYER metal4 ;
  RECT 2476.340 178.640 2477.460 179.760 ;
  LAYER metal3 ;
  RECT 2476.340 178.640 2477.460 179.760 ;
  LAYER metal2 ;
  RECT 2476.340 178.640 2477.460 179.760 ;
  LAYER metal1 ;
  RECT 2476.340 178.640 2477.460 179.760 ;
 END
END DIB88
PIN DOB88
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2462.700 178.640 2463.820 179.760 ;
  LAYER metal4 ;
  RECT 2462.700 178.640 2463.820 179.760 ;
  LAYER metal3 ;
  RECT 2462.700 178.640 2463.820 179.760 ;
  LAYER metal2 ;
  RECT 2462.700 178.640 2463.820 179.760 ;
  LAYER metal1 ;
  RECT 2462.700 178.640 2463.820 179.760 ;
 END
END DOB88
PIN DIB87
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2449.060 178.640 2450.180 179.760 ;
  LAYER metal4 ;
  RECT 2449.060 178.640 2450.180 179.760 ;
  LAYER metal3 ;
  RECT 2449.060 178.640 2450.180 179.760 ;
  LAYER metal2 ;
  RECT 2449.060 178.640 2450.180 179.760 ;
  LAYER metal1 ;
  RECT 2449.060 178.640 2450.180 179.760 ;
 END
END DIB87
PIN DOB87
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2436.040 178.640 2437.160 179.760 ;
  LAYER metal4 ;
  RECT 2436.040 178.640 2437.160 179.760 ;
  LAYER metal3 ;
  RECT 2436.040 178.640 2437.160 179.760 ;
  LAYER metal2 ;
  RECT 2436.040 178.640 2437.160 179.760 ;
  LAYER metal1 ;
  RECT 2436.040 178.640 2437.160 179.760 ;
 END
END DOB87
PIN DIB86
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2422.400 178.640 2423.520 179.760 ;
  LAYER metal4 ;
  RECT 2422.400 178.640 2423.520 179.760 ;
  LAYER metal3 ;
  RECT 2422.400 178.640 2423.520 179.760 ;
  LAYER metal2 ;
  RECT 2422.400 178.640 2423.520 179.760 ;
  LAYER metal1 ;
  RECT 2422.400 178.640 2423.520 179.760 ;
 END
END DIB86
PIN DOB86
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2408.760 178.640 2409.880 179.760 ;
  LAYER metal4 ;
  RECT 2408.760 178.640 2409.880 179.760 ;
  LAYER metal3 ;
  RECT 2408.760 178.640 2409.880 179.760 ;
  LAYER metal2 ;
  RECT 2408.760 178.640 2409.880 179.760 ;
  LAYER metal1 ;
  RECT 2408.760 178.640 2409.880 179.760 ;
 END
END DOB86
PIN DIB85
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2395.740 178.640 2396.860 179.760 ;
  LAYER metal4 ;
  RECT 2395.740 178.640 2396.860 179.760 ;
  LAYER metal3 ;
  RECT 2395.740 178.640 2396.860 179.760 ;
  LAYER metal2 ;
  RECT 2395.740 178.640 2396.860 179.760 ;
  LAYER metal1 ;
  RECT 2395.740 178.640 2396.860 179.760 ;
 END
END DIB85
PIN DOB85
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2382.100 178.640 2383.220 179.760 ;
  LAYER metal4 ;
  RECT 2382.100 178.640 2383.220 179.760 ;
  LAYER metal3 ;
  RECT 2382.100 178.640 2383.220 179.760 ;
  LAYER metal2 ;
  RECT 2382.100 178.640 2383.220 179.760 ;
  LAYER metal1 ;
  RECT 2382.100 178.640 2383.220 179.760 ;
 END
END DOB85
PIN DIB84
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2368.460 178.640 2369.580 179.760 ;
  LAYER metal4 ;
  RECT 2368.460 178.640 2369.580 179.760 ;
  LAYER metal3 ;
  RECT 2368.460 178.640 2369.580 179.760 ;
  LAYER metal2 ;
  RECT 2368.460 178.640 2369.580 179.760 ;
  LAYER metal1 ;
  RECT 2368.460 178.640 2369.580 179.760 ;
 END
END DIB84
PIN DOB84
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2355.440 178.640 2356.560 179.760 ;
  LAYER metal4 ;
  RECT 2355.440 178.640 2356.560 179.760 ;
  LAYER metal3 ;
  RECT 2355.440 178.640 2356.560 179.760 ;
  LAYER metal2 ;
  RECT 2355.440 178.640 2356.560 179.760 ;
  LAYER metal1 ;
  RECT 2355.440 178.640 2356.560 179.760 ;
 END
END DOB84
PIN DIB83
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2341.800 178.640 2342.920 179.760 ;
  LAYER metal4 ;
  RECT 2341.800 178.640 2342.920 179.760 ;
  LAYER metal3 ;
  RECT 2341.800 178.640 2342.920 179.760 ;
  LAYER metal2 ;
  RECT 2341.800 178.640 2342.920 179.760 ;
  LAYER metal1 ;
  RECT 2341.800 178.640 2342.920 179.760 ;
 END
END DIB83
PIN DOB83
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2328.160 178.640 2329.280 179.760 ;
  LAYER metal4 ;
  RECT 2328.160 178.640 2329.280 179.760 ;
  LAYER metal3 ;
  RECT 2328.160 178.640 2329.280 179.760 ;
  LAYER metal2 ;
  RECT 2328.160 178.640 2329.280 179.760 ;
  LAYER metal1 ;
  RECT 2328.160 178.640 2329.280 179.760 ;
 END
END DOB83
PIN DIB82
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2315.140 178.640 2316.260 179.760 ;
  LAYER metal4 ;
  RECT 2315.140 178.640 2316.260 179.760 ;
  LAYER metal3 ;
  RECT 2315.140 178.640 2316.260 179.760 ;
  LAYER metal2 ;
  RECT 2315.140 178.640 2316.260 179.760 ;
  LAYER metal1 ;
  RECT 2315.140 178.640 2316.260 179.760 ;
 END
END DIB82
PIN DOB82
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2301.500 178.640 2302.620 179.760 ;
  LAYER metal4 ;
  RECT 2301.500 178.640 2302.620 179.760 ;
  LAYER metal3 ;
  RECT 2301.500 178.640 2302.620 179.760 ;
  LAYER metal2 ;
  RECT 2301.500 178.640 2302.620 179.760 ;
  LAYER metal1 ;
  RECT 2301.500 178.640 2302.620 179.760 ;
 END
END DOB82
PIN DIB81
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2287.860 178.640 2288.980 179.760 ;
  LAYER metal4 ;
  RECT 2287.860 178.640 2288.980 179.760 ;
  LAYER metal3 ;
  RECT 2287.860 178.640 2288.980 179.760 ;
  LAYER metal2 ;
  RECT 2287.860 178.640 2288.980 179.760 ;
  LAYER metal1 ;
  RECT 2287.860 178.640 2288.980 179.760 ;
 END
END DIB81
PIN DOB81
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2274.840 178.640 2275.960 179.760 ;
  LAYER metal4 ;
  RECT 2274.840 178.640 2275.960 179.760 ;
  LAYER metal3 ;
  RECT 2274.840 178.640 2275.960 179.760 ;
  LAYER metal2 ;
  RECT 2274.840 178.640 2275.960 179.760 ;
  LAYER metal1 ;
  RECT 2274.840 178.640 2275.960 179.760 ;
 END
END DOB81
PIN DIB80
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2261.200 178.640 2262.320 179.760 ;
  LAYER metal4 ;
  RECT 2261.200 178.640 2262.320 179.760 ;
  LAYER metal3 ;
  RECT 2261.200 178.640 2262.320 179.760 ;
  LAYER metal2 ;
  RECT 2261.200 178.640 2262.320 179.760 ;
  LAYER metal1 ;
  RECT 2261.200 178.640 2262.320 179.760 ;
 END
END DIB80
PIN WEBN5
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2250.040 178.640 2251.160 179.760 ;
  LAYER metal4 ;
  RECT 2250.040 178.640 2251.160 179.760 ;
  LAYER metal3 ;
  RECT 2250.040 178.640 2251.160 179.760 ;
  LAYER metal2 ;
  RECT 2250.040 178.640 2251.160 179.760 ;
  LAYER metal1 ;
  RECT 2250.040 178.640 2251.160 179.760 ;
 END
END WEBN5
PIN DOB80
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2247.560 178.640 2248.680 179.760 ;
  LAYER metal4 ;
  RECT 2247.560 178.640 2248.680 179.760 ;
  LAYER metal3 ;
  RECT 2247.560 178.640 2248.680 179.760 ;
  LAYER metal2 ;
  RECT 2247.560 178.640 2248.680 179.760 ;
  LAYER metal1 ;
  RECT 2247.560 178.640 2248.680 179.760 ;
 END
END DOB80
PIN DIB79
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2234.540 178.640 2235.660 179.760 ;
  LAYER metal4 ;
  RECT 2234.540 178.640 2235.660 179.760 ;
  LAYER metal3 ;
  RECT 2234.540 178.640 2235.660 179.760 ;
  LAYER metal2 ;
  RECT 2234.540 178.640 2235.660 179.760 ;
  LAYER metal1 ;
  RECT 2234.540 178.640 2235.660 179.760 ;
 END
END DIB79
PIN DOB79
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2220.900 178.640 2222.020 179.760 ;
  LAYER metal4 ;
  RECT 2220.900 178.640 2222.020 179.760 ;
  LAYER metal3 ;
  RECT 2220.900 178.640 2222.020 179.760 ;
  LAYER metal2 ;
  RECT 2220.900 178.640 2222.020 179.760 ;
  LAYER metal1 ;
  RECT 2220.900 178.640 2222.020 179.760 ;
 END
END DOB79
PIN DIB78
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2207.260 178.640 2208.380 179.760 ;
  LAYER metal4 ;
  RECT 2207.260 178.640 2208.380 179.760 ;
  LAYER metal3 ;
  RECT 2207.260 178.640 2208.380 179.760 ;
  LAYER metal2 ;
  RECT 2207.260 178.640 2208.380 179.760 ;
  LAYER metal1 ;
  RECT 2207.260 178.640 2208.380 179.760 ;
 END
END DIB78
PIN DOB78
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2194.240 178.640 2195.360 179.760 ;
  LAYER metal4 ;
  RECT 2194.240 178.640 2195.360 179.760 ;
  LAYER metal3 ;
  RECT 2194.240 178.640 2195.360 179.760 ;
  LAYER metal2 ;
  RECT 2194.240 178.640 2195.360 179.760 ;
  LAYER metal1 ;
  RECT 2194.240 178.640 2195.360 179.760 ;
 END
END DOB78
PIN DIB77
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2180.600 178.640 2181.720 179.760 ;
  LAYER metal4 ;
  RECT 2180.600 178.640 2181.720 179.760 ;
  LAYER metal3 ;
  RECT 2180.600 178.640 2181.720 179.760 ;
  LAYER metal2 ;
  RECT 2180.600 178.640 2181.720 179.760 ;
  LAYER metal1 ;
  RECT 2180.600 178.640 2181.720 179.760 ;
 END
END DIB77
PIN DOB77
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2166.960 178.640 2168.080 179.760 ;
  LAYER metal4 ;
  RECT 2166.960 178.640 2168.080 179.760 ;
  LAYER metal3 ;
  RECT 2166.960 178.640 2168.080 179.760 ;
  LAYER metal2 ;
  RECT 2166.960 178.640 2168.080 179.760 ;
  LAYER metal1 ;
  RECT 2166.960 178.640 2168.080 179.760 ;
 END
END DOB77
PIN DIB76
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2153.940 178.640 2155.060 179.760 ;
  LAYER metal4 ;
  RECT 2153.940 178.640 2155.060 179.760 ;
  LAYER metal3 ;
  RECT 2153.940 178.640 2155.060 179.760 ;
  LAYER metal2 ;
  RECT 2153.940 178.640 2155.060 179.760 ;
  LAYER metal1 ;
  RECT 2153.940 178.640 2155.060 179.760 ;
 END
END DIB76
PIN DOB76
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2140.300 178.640 2141.420 179.760 ;
  LAYER metal4 ;
  RECT 2140.300 178.640 2141.420 179.760 ;
  LAYER metal3 ;
  RECT 2140.300 178.640 2141.420 179.760 ;
  LAYER metal2 ;
  RECT 2140.300 178.640 2141.420 179.760 ;
  LAYER metal1 ;
  RECT 2140.300 178.640 2141.420 179.760 ;
 END
END DOB76
PIN DIB75
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2126.660 178.640 2127.780 179.760 ;
  LAYER metal4 ;
  RECT 2126.660 178.640 2127.780 179.760 ;
  LAYER metal3 ;
  RECT 2126.660 178.640 2127.780 179.760 ;
  LAYER metal2 ;
  RECT 2126.660 178.640 2127.780 179.760 ;
  LAYER metal1 ;
  RECT 2126.660 178.640 2127.780 179.760 ;
 END
END DIB75
PIN DOB75
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2113.640 178.640 2114.760 179.760 ;
  LAYER metal4 ;
  RECT 2113.640 178.640 2114.760 179.760 ;
  LAYER metal3 ;
  RECT 2113.640 178.640 2114.760 179.760 ;
  LAYER metal2 ;
  RECT 2113.640 178.640 2114.760 179.760 ;
  LAYER metal1 ;
  RECT 2113.640 178.640 2114.760 179.760 ;
 END
END DOB75
PIN DIB74
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2100.000 178.640 2101.120 179.760 ;
  LAYER metal4 ;
  RECT 2100.000 178.640 2101.120 179.760 ;
  LAYER metal3 ;
  RECT 2100.000 178.640 2101.120 179.760 ;
  LAYER metal2 ;
  RECT 2100.000 178.640 2101.120 179.760 ;
  LAYER metal1 ;
  RECT 2100.000 178.640 2101.120 179.760 ;
 END
END DIB74
PIN DOB74
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2086.360 178.640 2087.480 179.760 ;
  LAYER metal4 ;
  RECT 2086.360 178.640 2087.480 179.760 ;
  LAYER metal3 ;
  RECT 2086.360 178.640 2087.480 179.760 ;
  LAYER metal2 ;
  RECT 2086.360 178.640 2087.480 179.760 ;
  LAYER metal1 ;
  RECT 2086.360 178.640 2087.480 179.760 ;
 END
END DOB74
PIN DIB73
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2072.720 178.640 2073.840 179.760 ;
  LAYER metal4 ;
  RECT 2072.720 178.640 2073.840 179.760 ;
  LAYER metal3 ;
  RECT 2072.720 178.640 2073.840 179.760 ;
  LAYER metal2 ;
  RECT 2072.720 178.640 2073.840 179.760 ;
  LAYER metal1 ;
  RECT 2072.720 178.640 2073.840 179.760 ;
 END
END DIB73
PIN DOB73
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2059.700 178.640 2060.820 179.760 ;
  LAYER metal4 ;
  RECT 2059.700 178.640 2060.820 179.760 ;
  LAYER metal3 ;
  RECT 2059.700 178.640 2060.820 179.760 ;
  LAYER metal2 ;
  RECT 2059.700 178.640 2060.820 179.760 ;
  LAYER metal1 ;
  RECT 2059.700 178.640 2060.820 179.760 ;
 END
END DOB73
PIN DIB72
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2046.060 178.640 2047.180 179.760 ;
  LAYER metal4 ;
  RECT 2046.060 178.640 2047.180 179.760 ;
  LAYER metal3 ;
  RECT 2046.060 178.640 2047.180 179.760 ;
  LAYER metal2 ;
  RECT 2046.060 178.640 2047.180 179.760 ;
  LAYER metal1 ;
  RECT 2046.060 178.640 2047.180 179.760 ;
 END
END DIB72
PIN DOB72
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2032.420 178.640 2033.540 179.760 ;
  LAYER metal4 ;
  RECT 2032.420 178.640 2033.540 179.760 ;
  LAYER metal3 ;
  RECT 2032.420 178.640 2033.540 179.760 ;
  LAYER metal2 ;
  RECT 2032.420 178.640 2033.540 179.760 ;
  LAYER metal1 ;
  RECT 2032.420 178.640 2033.540 179.760 ;
 END
END DOB72
PIN DIB71
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2019.400 178.640 2020.520 179.760 ;
  LAYER metal4 ;
  RECT 2019.400 178.640 2020.520 179.760 ;
  LAYER metal3 ;
  RECT 2019.400 178.640 2020.520 179.760 ;
  LAYER metal2 ;
  RECT 2019.400 178.640 2020.520 179.760 ;
  LAYER metal1 ;
  RECT 2019.400 178.640 2020.520 179.760 ;
 END
END DIB71
PIN DOB71
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2005.760 178.640 2006.880 179.760 ;
  LAYER metal4 ;
  RECT 2005.760 178.640 2006.880 179.760 ;
  LAYER metal3 ;
  RECT 2005.760 178.640 2006.880 179.760 ;
  LAYER metal2 ;
  RECT 2005.760 178.640 2006.880 179.760 ;
  LAYER metal1 ;
  RECT 2005.760 178.640 2006.880 179.760 ;
 END
END DOB71
PIN DIB70
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1992.120 178.640 1993.240 179.760 ;
  LAYER metal4 ;
  RECT 1992.120 178.640 1993.240 179.760 ;
  LAYER metal3 ;
  RECT 1992.120 178.640 1993.240 179.760 ;
  LAYER metal2 ;
  RECT 1992.120 178.640 1993.240 179.760 ;
  LAYER metal1 ;
  RECT 1992.120 178.640 1993.240 179.760 ;
 END
END DIB70
PIN DOB70
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1979.100 178.640 1980.220 179.760 ;
  LAYER metal4 ;
  RECT 1979.100 178.640 1980.220 179.760 ;
  LAYER metal3 ;
  RECT 1979.100 178.640 1980.220 179.760 ;
  LAYER metal2 ;
  RECT 1979.100 178.640 1980.220 179.760 ;
  LAYER metal1 ;
  RECT 1979.100 178.640 1980.220 179.760 ;
 END
END DOB70
PIN DIB69
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1965.460 178.640 1966.580 179.760 ;
  LAYER metal4 ;
  RECT 1965.460 178.640 1966.580 179.760 ;
  LAYER metal3 ;
  RECT 1965.460 178.640 1966.580 179.760 ;
  LAYER metal2 ;
  RECT 1965.460 178.640 1966.580 179.760 ;
  LAYER metal1 ;
  RECT 1965.460 178.640 1966.580 179.760 ;
 END
END DIB69
PIN DOB69
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1951.820 178.640 1952.940 179.760 ;
  LAYER metal4 ;
  RECT 1951.820 178.640 1952.940 179.760 ;
  LAYER metal3 ;
  RECT 1951.820 178.640 1952.940 179.760 ;
  LAYER metal2 ;
  RECT 1951.820 178.640 1952.940 179.760 ;
  LAYER metal1 ;
  RECT 1951.820 178.640 1952.940 179.760 ;
 END
END DOB69
PIN DIB68
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1938.800 178.640 1939.920 179.760 ;
  LAYER metal4 ;
  RECT 1938.800 178.640 1939.920 179.760 ;
  LAYER metal3 ;
  RECT 1938.800 178.640 1939.920 179.760 ;
  LAYER metal2 ;
  RECT 1938.800 178.640 1939.920 179.760 ;
  LAYER metal1 ;
  RECT 1938.800 178.640 1939.920 179.760 ;
 END
END DIB68
PIN DOB68
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1925.160 178.640 1926.280 179.760 ;
  LAYER metal4 ;
  RECT 1925.160 178.640 1926.280 179.760 ;
  LAYER metal3 ;
  RECT 1925.160 178.640 1926.280 179.760 ;
  LAYER metal2 ;
  RECT 1925.160 178.640 1926.280 179.760 ;
  LAYER metal1 ;
  RECT 1925.160 178.640 1926.280 179.760 ;
 END
END DOB68
PIN DIB67
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1911.520 178.640 1912.640 179.760 ;
  LAYER metal4 ;
  RECT 1911.520 178.640 1912.640 179.760 ;
  LAYER metal3 ;
  RECT 1911.520 178.640 1912.640 179.760 ;
  LAYER metal2 ;
  RECT 1911.520 178.640 1912.640 179.760 ;
  LAYER metal1 ;
  RECT 1911.520 178.640 1912.640 179.760 ;
 END
END DIB67
PIN DOB67
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1898.500 178.640 1899.620 179.760 ;
  LAYER metal4 ;
  RECT 1898.500 178.640 1899.620 179.760 ;
  LAYER metal3 ;
  RECT 1898.500 178.640 1899.620 179.760 ;
  LAYER metal2 ;
  RECT 1898.500 178.640 1899.620 179.760 ;
  LAYER metal1 ;
  RECT 1898.500 178.640 1899.620 179.760 ;
 END
END DOB67
PIN DIB66
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1884.860 178.640 1885.980 179.760 ;
  LAYER metal4 ;
  RECT 1884.860 178.640 1885.980 179.760 ;
  LAYER metal3 ;
  RECT 1884.860 178.640 1885.980 179.760 ;
  LAYER metal2 ;
  RECT 1884.860 178.640 1885.980 179.760 ;
  LAYER metal1 ;
  RECT 1884.860 178.640 1885.980 179.760 ;
 END
END DIB66
PIN DOB66
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1871.220 178.640 1872.340 179.760 ;
  LAYER metal4 ;
  RECT 1871.220 178.640 1872.340 179.760 ;
  LAYER metal3 ;
  RECT 1871.220 178.640 1872.340 179.760 ;
  LAYER metal2 ;
  RECT 1871.220 178.640 1872.340 179.760 ;
  LAYER metal1 ;
  RECT 1871.220 178.640 1872.340 179.760 ;
 END
END DOB66
PIN DIB65
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1858.200 178.640 1859.320 179.760 ;
  LAYER metal4 ;
  RECT 1858.200 178.640 1859.320 179.760 ;
  LAYER metal3 ;
  RECT 1858.200 178.640 1859.320 179.760 ;
  LAYER metal2 ;
  RECT 1858.200 178.640 1859.320 179.760 ;
  LAYER metal1 ;
  RECT 1858.200 178.640 1859.320 179.760 ;
 END
END DIB65
PIN DOB65
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1844.560 178.640 1845.680 179.760 ;
  LAYER metal4 ;
  RECT 1844.560 178.640 1845.680 179.760 ;
  LAYER metal3 ;
  RECT 1844.560 178.640 1845.680 179.760 ;
  LAYER metal2 ;
  RECT 1844.560 178.640 1845.680 179.760 ;
  LAYER metal1 ;
  RECT 1844.560 178.640 1845.680 179.760 ;
 END
END DOB65
PIN DIB64
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1830.920 178.640 1832.040 179.760 ;
  LAYER metal4 ;
  RECT 1830.920 178.640 1832.040 179.760 ;
  LAYER metal3 ;
  RECT 1830.920 178.640 1832.040 179.760 ;
  LAYER metal2 ;
  RECT 1830.920 178.640 1832.040 179.760 ;
  LAYER metal1 ;
  RECT 1830.920 178.640 1832.040 179.760 ;
 END
END DIB64
PIN WEBN4
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1819.760 178.640 1820.880 179.760 ;
  LAYER metal4 ;
  RECT 1819.760 178.640 1820.880 179.760 ;
  LAYER metal3 ;
  RECT 1819.760 178.640 1820.880 179.760 ;
  LAYER metal2 ;
  RECT 1819.760 178.640 1820.880 179.760 ;
  LAYER metal1 ;
  RECT 1819.760 178.640 1820.880 179.760 ;
 END
END WEBN4
PIN DOB64
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1817.900 178.640 1819.020 179.760 ;
  LAYER metal4 ;
  RECT 1817.900 178.640 1819.020 179.760 ;
  LAYER metal3 ;
  RECT 1817.900 178.640 1819.020 179.760 ;
  LAYER metal2 ;
  RECT 1817.900 178.640 1819.020 179.760 ;
  LAYER metal1 ;
  RECT 1817.900 178.640 1819.020 179.760 ;
 END
END DOB64
PIN OEB
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1790.620 178.640 1791.740 179.760 ;
  LAYER metal4 ;
  RECT 1790.620 178.640 1791.740 179.760 ;
  LAYER metal3 ;
  RECT 1790.620 178.640 1791.740 179.760 ;
  LAYER metal2 ;
  RECT 1790.620 178.640 1791.740 179.760 ;
  LAYER metal1 ;
  RECT 1790.620 178.640 1791.740 179.760 ;
 END
END OEB
PIN CKB
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1777.600 178.640 1778.720 179.760 ;
  LAYER metal4 ;
  RECT 1777.600 178.640 1778.720 179.760 ;
  LAYER metal3 ;
  RECT 1777.600 178.640 1778.720 179.760 ;
  LAYER metal2 ;
  RECT 1777.600 178.640 1778.720 179.760 ;
  LAYER metal1 ;
  RECT 1777.600 178.640 1778.720 179.760 ;
 END
END CKB
PIN CSB
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1775.740 178.640 1776.860 179.760 ;
  LAYER metal4 ;
  RECT 1775.740 178.640 1776.860 179.760 ;
  LAYER metal3 ;
  RECT 1775.740 178.640 1776.860 179.760 ;
  LAYER metal2 ;
  RECT 1775.740 178.640 1776.860 179.760 ;
  LAYER metal1 ;
  RECT 1775.740 178.640 1776.860 179.760 ;
 END
END CSB
PIN B2
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1768.920 178.640 1770.040 179.760 ;
  LAYER metal4 ;
  RECT 1768.920 178.640 1770.040 179.760 ;
  LAYER metal3 ;
  RECT 1768.920 178.640 1770.040 179.760 ;
  LAYER metal2 ;
  RECT 1768.920 178.640 1770.040 179.760 ;
  LAYER metal1 ;
  RECT 1768.920 178.640 1770.040 179.760 ;
 END
END B2
PIN B1
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1763.960 178.640 1765.080 179.760 ;
  LAYER metal4 ;
  RECT 1763.960 178.640 1765.080 179.760 ;
  LAYER metal3 ;
  RECT 1763.960 178.640 1765.080 179.760 ;
  LAYER metal2 ;
  RECT 1763.960 178.640 1765.080 179.760 ;
  LAYER metal1 ;
  RECT 1763.960 178.640 1765.080 179.760 ;
 END
END B1
PIN B0
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1761.480 178.640 1762.600 179.760 ;
  LAYER metal4 ;
  RECT 1761.480 178.640 1762.600 179.760 ;
  LAYER metal3 ;
  RECT 1761.480 178.640 1762.600 179.760 ;
  LAYER metal2 ;
  RECT 1761.480 178.640 1762.600 179.760 ;
  LAYER metal1 ;
  RECT 1761.480 178.640 1762.600 179.760 ;
 END
END B0
PIN B5
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1753.420 178.640 1754.540 179.760 ;
  LAYER metal4 ;
  RECT 1753.420 178.640 1754.540 179.760 ;
  LAYER metal3 ;
  RECT 1753.420 178.640 1754.540 179.760 ;
  LAYER metal2 ;
  RECT 1753.420 178.640 1754.540 179.760 ;
  LAYER metal1 ;
  RECT 1753.420 178.640 1754.540 179.760 ;
 END
END B5
PIN B4
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1747.840 178.640 1748.960 179.760 ;
  LAYER metal4 ;
  RECT 1747.840 178.640 1748.960 179.760 ;
  LAYER metal3 ;
  RECT 1747.840 178.640 1748.960 179.760 ;
  LAYER metal2 ;
  RECT 1747.840 178.640 1748.960 179.760 ;
  LAYER metal1 ;
  RECT 1747.840 178.640 1748.960 179.760 ;
 END
END B4
PIN B3
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1741.640 178.640 1742.760 179.760 ;
  LAYER metal4 ;
  RECT 1741.640 178.640 1742.760 179.760 ;
  LAYER metal3 ;
  RECT 1741.640 178.640 1742.760 179.760 ;
  LAYER metal2 ;
  RECT 1741.640 178.640 1742.760 179.760 ;
  LAYER metal1 ;
  RECT 1741.640 178.640 1742.760 179.760 ;
 END
END B3
PIN DIB63
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1719.320 178.640 1720.440 179.760 ;
  LAYER metal4 ;
  RECT 1719.320 178.640 1720.440 179.760 ;
  LAYER metal3 ;
  RECT 1719.320 178.640 1720.440 179.760 ;
  LAYER metal2 ;
  RECT 1719.320 178.640 1720.440 179.760 ;
  LAYER metal1 ;
  RECT 1719.320 178.640 1720.440 179.760 ;
 END
END DIB63
PIN DOB63
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1706.300 178.640 1707.420 179.760 ;
  LAYER metal4 ;
  RECT 1706.300 178.640 1707.420 179.760 ;
  LAYER metal3 ;
  RECT 1706.300 178.640 1707.420 179.760 ;
  LAYER metal2 ;
  RECT 1706.300 178.640 1707.420 179.760 ;
  LAYER metal1 ;
  RECT 1706.300 178.640 1707.420 179.760 ;
 END
END DOB63
PIN DIB62
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1692.660 178.640 1693.780 179.760 ;
  LAYER metal4 ;
  RECT 1692.660 178.640 1693.780 179.760 ;
  LAYER metal3 ;
  RECT 1692.660 178.640 1693.780 179.760 ;
  LAYER metal2 ;
  RECT 1692.660 178.640 1693.780 179.760 ;
  LAYER metal1 ;
  RECT 1692.660 178.640 1693.780 179.760 ;
 END
END DIB62
PIN DOB62
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1679.020 178.640 1680.140 179.760 ;
  LAYER metal4 ;
  RECT 1679.020 178.640 1680.140 179.760 ;
  LAYER metal3 ;
  RECT 1679.020 178.640 1680.140 179.760 ;
  LAYER metal2 ;
  RECT 1679.020 178.640 1680.140 179.760 ;
  LAYER metal1 ;
  RECT 1679.020 178.640 1680.140 179.760 ;
 END
END DOB62
PIN DIB61
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1666.000 178.640 1667.120 179.760 ;
  LAYER metal4 ;
  RECT 1666.000 178.640 1667.120 179.760 ;
  LAYER metal3 ;
  RECT 1666.000 178.640 1667.120 179.760 ;
  LAYER metal2 ;
  RECT 1666.000 178.640 1667.120 179.760 ;
  LAYER metal1 ;
  RECT 1666.000 178.640 1667.120 179.760 ;
 END
END DIB61
PIN DOB61
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1652.360 178.640 1653.480 179.760 ;
  LAYER metal4 ;
  RECT 1652.360 178.640 1653.480 179.760 ;
  LAYER metal3 ;
  RECT 1652.360 178.640 1653.480 179.760 ;
  LAYER metal2 ;
  RECT 1652.360 178.640 1653.480 179.760 ;
  LAYER metal1 ;
  RECT 1652.360 178.640 1653.480 179.760 ;
 END
END DOB61
PIN DIB60
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1638.720 178.640 1639.840 179.760 ;
  LAYER metal4 ;
  RECT 1638.720 178.640 1639.840 179.760 ;
  LAYER metal3 ;
  RECT 1638.720 178.640 1639.840 179.760 ;
  LAYER metal2 ;
  RECT 1638.720 178.640 1639.840 179.760 ;
  LAYER metal1 ;
  RECT 1638.720 178.640 1639.840 179.760 ;
 END
END DIB60
PIN DOB60
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1625.700 178.640 1626.820 179.760 ;
  LAYER metal4 ;
  RECT 1625.700 178.640 1626.820 179.760 ;
  LAYER metal3 ;
  RECT 1625.700 178.640 1626.820 179.760 ;
  LAYER metal2 ;
  RECT 1625.700 178.640 1626.820 179.760 ;
  LAYER metal1 ;
  RECT 1625.700 178.640 1626.820 179.760 ;
 END
END DOB60
PIN DIB59
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1612.060 178.640 1613.180 179.760 ;
  LAYER metal4 ;
  RECT 1612.060 178.640 1613.180 179.760 ;
  LAYER metal3 ;
  RECT 1612.060 178.640 1613.180 179.760 ;
  LAYER metal2 ;
  RECT 1612.060 178.640 1613.180 179.760 ;
  LAYER metal1 ;
  RECT 1612.060 178.640 1613.180 179.760 ;
 END
END DIB59
PIN DOB59
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1598.420 178.640 1599.540 179.760 ;
  LAYER metal4 ;
  RECT 1598.420 178.640 1599.540 179.760 ;
  LAYER metal3 ;
  RECT 1598.420 178.640 1599.540 179.760 ;
  LAYER metal2 ;
  RECT 1598.420 178.640 1599.540 179.760 ;
  LAYER metal1 ;
  RECT 1598.420 178.640 1599.540 179.760 ;
 END
END DOB59
PIN DIB58
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1585.400 178.640 1586.520 179.760 ;
  LAYER metal4 ;
  RECT 1585.400 178.640 1586.520 179.760 ;
  LAYER metal3 ;
  RECT 1585.400 178.640 1586.520 179.760 ;
  LAYER metal2 ;
  RECT 1585.400 178.640 1586.520 179.760 ;
  LAYER metal1 ;
  RECT 1585.400 178.640 1586.520 179.760 ;
 END
END DIB58
PIN DOB58
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1571.760 178.640 1572.880 179.760 ;
  LAYER metal4 ;
  RECT 1571.760 178.640 1572.880 179.760 ;
  LAYER metal3 ;
  RECT 1571.760 178.640 1572.880 179.760 ;
  LAYER metal2 ;
  RECT 1571.760 178.640 1572.880 179.760 ;
  LAYER metal1 ;
  RECT 1571.760 178.640 1572.880 179.760 ;
 END
END DOB58
PIN DIB57
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1558.120 178.640 1559.240 179.760 ;
  LAYER metal4 ;
  RECT 1558.120 178.640 1559.240 179.760 ;
  LAYER metal3 ;
  RECT 1558.120 178.640 1559.240 179.760 ;
  LAYER metal2 ;
  RECT 1558.120 178.640 1559.240 179.760 ;
  LAYER metal1 ;
  RECT 1558.120 178.640 1559.240 179.760 ;
 END
END DIB57
PIN DOB57
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1545.100 178.640 1546.220 179.760 ;
  LAYER metal4 ;
  RECT 1545.100 178.640 1546.220 179.760 ;
  LAYER metal3 ;
  RECT 1545.100 178.640 1546.220 179.760 ;
  LAYER metal2 ;
  RECT 1545.100 178.640 1546.220 179.760 ;
  LAYER metal1 ;
  RECT 1545.100 178.640 1546.220 179.760 ;
 END
END DOB57
PIN DIB56
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1531.460 178.640 1532.580 179.760 ;
  LAYER metal4 ;
  RECT 1531.460 178.640 1532.580 179.760 ;
  LAYER metal3 ;
  RECT 1531.460 178.640 1532.580 179.760 ;
  LAYER metal2 ;
  RECT 1531.460 178.640 1532.580 179.760 ;
  LAYER metal1 ;
  RECT 1531.460 178.640 1532.580 179.760 ;
 END
END DIB56
PIN DOB56
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1517.820 178.640 1518.940 179.760 ;
  LAYER metal4 ;
  RECT 1517.820 178.640 1518.940 179.760 ;
  LAYER metal3 ;
  RECT 1517.820 178.640 1518.940 179.760 ;
  LAYER metal2 ;
  RECT 1517.820 178.640 1518.940 179.760 ;
  LAYER metal1 ;
  RECT 1517.820 178.640 1518.940 179.760 ;
 END
END DOB56
PIN DIB55
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1504.800 178.640 1505.920 179.760 ;
  LAYER metal4 ;
  RECT 1504.800 178.640 1505.920 179.760 ;
  LAYER metal3 ;
  RECT 1504.800 178.640 1505.920 179.760 ;
  LAYER metal2 ;
  RECT 1504.800 178.640 1505.920 179.760 ;
  LAYER metal1 ;
  RECT 1504.800 178.640 1505.920 179.760 ;
 END
END DIB55
PIN DOB55
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1491.160 178.640 1492.280 179.760 ;
  LAYER metal4 ;
  RECT 1491.160 178.640 1492.280 179.760 ;
  LAYER metal3 ;
  RECT 1491.160 178.640 1492.280 179.760 ;
  LAYER metal2 ;
  RECT 1491.160 178.640 1492.280 179.760 ;
  LAYER metal1 ;
  RECT 1491.160 178.640 1492.280 179.760 ;
 END
END DOB55
PIN DIB54
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1477.520 178.640 1478.640 179.760 ;
  LAYER metal4 ;
  RECT 1477.520 178.640 1478.640 179.760 ;
  LAYER metal3 ;
  RECT 1477.520 178.640 1478.640 179.760 ;
  LAYER metal2 ;
  RECT 1477.520 178.640 1478.640 179.760 ;
  LAYER metal1 ;
  RECT 1477.520 178.640 1478.640 179.760 ;
 END
END DIB54
PIN DOB54
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1464.500 178.640 1465.620 179.760 ;
  LAYER metal4 ;
  RECT 1464.500 178.640 1465.620 179.760 ;
  LAYER metal3 ;
  RECT 1464.500 178.640 1465.620 179.760 ;
  LAYER metal2 ;
  RECT 1464.500 178.640 1465.620 179.760 ;
  LAYER metal1 ;
  RECT 1464.500 178.640 1465.620 179.760 ;
 END
END DOB54
PIN DIB53
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1450.860 178.640 1451.980 179.760 ;
  LAYER metal4 ;
  RECT 1450.860 178.640 1451.980 179.760 ;
  LAYER metal3 ;
  RECT 1450.860 178.640 1451.980 179.760 ;
  LAYER metal2 ;
  RECT 1450.860 178.640 1451.980 179.760 ;
  LAYER metal1 ;
  RECT 1450.860 178.640 1451.980 179.760 ;
 END
END DIB53
PIN DOB53
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1437.220 178.640 1438.340 179.760 ;
  LAYER metal4 ;
  RECT 1437.220 178.640 1438.340 179.760 ;
  LAYER metal3 ;
  RECT 1437.220 178.640 1438.340 179.760 ;
  LAYER metal2 ;
  RECT 1437.220 178.640 1438.340 179.760 ;
  LAYER metal1 ;
  RECT 1437.220 178.640 1438.340 179.760 ;
 END
END DOB53
PIN DIB52
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1424.200 178.640 1425.320 179.760 ;
  LAYER metal4 ;
  RECT 1424.200 178.640 1425.320 179.760 ;
  LAYER metal3 ;
  RECT 1424.200 178.640 1425.320 179.760 ;
  LAYER metal2 ;
  RECT 1424.200 178.640 1425.320 179.760 ;
  LAYER metal1 ;
  RECT 1424.200 178.640 1425.320 179.760 ;
 END
END DIB52
PIN DOB52
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1410.560 178.640 1411.680 179.760 ;
  LAYER metal4 ;
  RECT 1410.560 178.640 1411.680 179.760 ;
  LAYER metal3 ;
  RECT 1410.560 178.640 1411.680 179.760 ;
  LAYER metal2 ;
  RECT 1410.560 178.640 1411.680 179.760 ;
  LAYER metal1 ;
  RECT 1410.560 178.640 1411.680 179.760 ;
 END
END DOB52
PIN DIB51
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1396.920 178.640 1398.040 179.760 ;
  LAYER metal4 ;
  RECT 1396.920 178.640 1398.040 179.760 ;
  LAYER metal3 ;
  RECT 1396.920 178.640 1398.040 179.760 ;
  LAYER metal2 ;
  RECT 1396.920 178.640 1398.040 179.760 ;
  LAYER metal1 ;
  RECT 1396.920 178.640 1398.040 179.760 ;
 END
END DIB51
PIN DOB51
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1383.900 178.640 1385.020 179.760 ;
  LAYER metal4 ;
  RECT 1383.900 178.640 1385.020 179.760 ;
  LAYER metal3 ;
  RECT 1383.900 178.640 1385.020 179.760 ;
  LAYER metal2 ;
  RECT 1383.900 178.640 1385.020 179.760 ;
  LAYER metal1 ;
  RECT 1383.900 178.640 1385.020 179.760 ;
 END
END DOB51
PIN DIB50
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1370.260 178.640 1371.380 179.760 ;
  LAYER metal4 ;
  RECT 1370.260 178.640 1371.380 179.760 ;
  LAYER metal3 ;
  RECT 1370.260 178.640 1371.380 179.760 ;
  LAYER metal2 ;
  RECT 1370.260 178.640 1371.380 179.760 ;
  LAYER metal1 ;
  RECT 1370.260 178.640 1371.380 179.760 ;
 END
END DIB50
PIN DOB50
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1356.620 178.640 1357.740 179.760 ;
  LAYER metal4 ;
  RECT 1356.620 178.640 1357.740 179.760 ;
  LAYER metal3 ;
  RECT 1356.620 178.640 1357.740 179.760 ;
  LAYER metal2 ;
  RECT 1356.620 178.640 1357.740 179.760 ;
  LAYER metal1 ;
  RECT 1356.620 178.640 1357.740 179.760 ;
 END
END DOB50
PIN DIB49
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1343.600 178.640 1344.720 179.760 ;
  LAYER metal4 ;
  RECT 1343.600 178.640 1344.720 179.760 ;
  LAYER metal3 ;
  RECT 1343.600 178.640 1344.720 179.760 ;
  LAYER metal2 ;
  RECT 1343.600 178.640 1344.720 179.760 ;
  LAYER metal1 ;
  RECT 1343.600 178.640 1344.720 179.760 ;
 END
END DIB49
PIN DOB49
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1329.960 178.640 1331.080 179.760 ;
  LAYER metal4 ;
  RECT 1329.960 178.640 1331.080 179.760 ;
  LAYER metal3 ;
  RECT 1329.960 178.640 1331.080 179.760 ;
  LAYER metal2 ;
  RECT 1329.960 178.640 1331.080 179.760 ;
  LAYER metal1 ;
  RECT 1329.960 178.640 1331.080 179.760 ;
 END
END DOB49
PIN DIB48
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1316.320 178.640 1317.440 179.760 ;
  LAYER metal4 ;
  RECT 1316.320 178.640 1317.440 179.760 ;
  LAYER metal3 ;
  RECT 1316.320 178.640 1317.440 179.760 ;
  LAYER metal2 ;
  RECT 1316.320 178.640 1317.440 179.760 ;
  LAYER metal1 ;
  RECT 1316.320 178.640 1317.440 179.760 ;
 END
END DIB48
PIN WEBN3
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1305.160 178.640 1306.280 179.760 ;
  LAYER metal4 ;
  RECT 1305.160 178.640 1306.280 179.760 ;
  LAYER metal3 ;
  RECT 1305.160 178.640 1306.280 179.760 ;
  LAYER metal2 ;
  RECT 1305.160 178.640 1306.280 179.760 ;
  LAYER metal1 ;
  RECT 1305.160 178.640 1306.280 179.760 ;
 END
END WEBN3
PIN DOB48
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1302.680 178.640 1303.800 179.760 ;
  LAYER metal4 ;
  RECT 1302.680 178.640 1303.800 179.760 ;
  LAYER metal3 ;
  RECT 1302.680 178.640 1303.800 179.760 ;
  LAYER metal2 ;
  RECT 1302.680 178.640 1303.800 179.760 ;
  LAYER metal1 ;
  RECT 1302.680 178.640 1303.800 179.760 ;
 END
END DOB48
PIN DIB47
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1289.660 178.640 1290.780 179.760 ;
  LAYER metal4 ;
  RECT 1289.660 178.640 1290.780 179.760 ;
  LAYER metal3 ;
  RECT 1289.660 178.640 1290.780 179.760 ;
  LAYER metal2 ;
  RECT 1289.660 178.640 1290.780 179.760 ;
  LAYER metal1 ;
  RECT 1289.660 178.640 1290.780 179.760 ;
 END
END DIB47
PIN DOB47
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1276.020 178.640 1277.140 179.760 ;
  LAYER metal4 ;
  RECT 1276.020 178.640 1277.140 179.760 ;
  LAYER metal3 ;
  RECT 1276.020 178.640 1277.140 179.760 ;
  LAYER metal2 ;
  RECT 1276.020 178.640 1277.140 179.760 ;
  LAYER metal1 ;
  RECT 1276.020 178.640 1277.140 179.760 ;
 END
END DOB47
PIN DIB46
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1262.380 178.640 1263.500 179.760 ;
  LAYER metal4 ;
  RECT 1262.380 178.640 1263.500 179.760 ;
  LAYER metal3 ;
  RECT 1262.380 178.640 1263.500 179.760 ;
  LAYER metal2 ;
  RECT 1262.380 178.640 1263.500 179.760 ;
  LAYER metal1 ;
  RECT 1262.380 178.640 1263.500 179.760 ;
 END
END DIB46
PIN DOB46
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1249.360 178.640 1250.480 179.760 ;
  LAYER metal4 ;
  RECT 1249.360 178.640 1250.480 179.760 ;
  LAYER metal3 ;
  RECT 1249.360 178.640 1250.480 179.760 ;
  LAYER metal2 ;
  RECT 1249.360 178.640 1250.480 179.760 ;
  LAYER metal1 ;
  RECT 1249.360 178.640 1250.480 179.760 ;
 END
END DOB46
PIN DIB45
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1235.720 178.640 1236.840 179.760 ;
  LAYER metal4 ;
  RECT 1235.720 178.640 1236.840 179.760 ;
  LAYER metal3 ;
  RECT 1235.720 178.640 1236.840 179.760 ;
  LAYER metal2 ;
  RECT 1235.720 178.640 1236.840 179.760 ;
  LAYER metal1 ;
  RECT 1235.720 178.640 1236.840 179.760 ;
 END
END DIB45
PIN DOB45
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1222.080 178.640 1223.200 179.760 ;
  LAYER metal4 ;
  RECT 1222.080 178.640 1223.200 179.760 ;
  LAYER metal3 ;
  RECT 1222.080 178.640 1223.200 179.760 ;
  LAYER metal2 ;
  RECT 1222.080 178.640 1223.200 179.760 ;
  LAYER metal1 ;
  RECT 1222.080 178.640 1223.200 179.760 ;
 END
END DOB45
PIN DIB44
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1209.060 178.640 1210.180 179.760 ;
  LAYER metal4 ;
  RECT 1209.060 178.640 1210.180 179.760 ;
  LAYER metal3 ;
  RECT 1209.060 178.640 1210.180 179.760 ;
  LAYER metal2 ;
  RECT 1209.060 178.640 1210.180 179.760 ;
  LAYER metal1 ;
  RECT 1209.060 178.640 1210.180 179.760 ;
 END
END DIB44
PIN DOB44
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1195.420 178.640 1196.540 179.760 ;
  LAYER metal4 ;
  RECT 1195.420 178.640 1196.540 179.760 ;
  LAYER metal3 ;
  RECT 1195.420 178.640 1196.540 179.760 ;
  LAYER metal2 ;
  RECT 1195.420 178.640 1196.540 179.760 ;
  LAYER metal1 ;
  RECT 1195.420 178.640 1196.540 179.760 ;
 END
END DOB44
PIN DIB43
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1181.780 178.640 1182.900 179.760 ;
  LAYER metal4 ;
  RECT 1181.780 178.640 1182.900 179.760 ;
  LAYER metal3 ;
  RECT 1181.780 178.640 1182.900 179.760 ;
  LAYER metal2 ;
  RECT 1181.780 178.640 1182.900 179.760 ;
  LAYER metal1 ;
  RECT 1181.780 178.640 1182.900 179.760 ;
 END
END DIB43
PIN DOB43
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1168.760 178.640 1169.880 179.760 ;
  LAYER metal4 ;
  RECT 1168.760 178.640 1169.880 179.760 ;
  LAYER metal3 ;
  RECT 1168.760 178.640 1169.880 179.760 ;
  LAYER metal2 ;
  RECT 1168.760 178.640 1169.880 179.760 ;
  LAYER metal1 ;
  RECT 1168.760 178.640 1169.880 179.760 ;
 END
END DOB43
PIN DIB42
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1155.120 178.640 1156.240 179.760 ;
  LAYER metal4 ;
  RECT 1155.120 178.640 1156.240 179.760 ;
  LAYER metal3 ;
  RECT 1155.120 178.640 1156.240 179.760 ;
  LAYER metal2 ;
  RECT 1155.120 178.640 1156.240 179.760 ;
  LAYER metal1 ;
  RECT 1155.120 178.640 1156.240 179.760 ;
 END
END DIB42
PIN DOB42
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1141.480 178.640 1142.600 179.760 ;
  LAYER metal4 ;
  RECT 1141.480 178.640 1142.600 179.760 ;
  LAYER metal3 ;
  RECT 1141.480 178.640 1142.600 179.760 ;
  LAYER metal2 ;
  RECT 1141.480 178.640 1142.600 179.760 ;
  LAYER metal1 ;
  RECT 1141.480 178.640 1142.600 179.760 ;
 END
END DOB42
PIN DIB41
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1128.460 178.640 1129.580 179.760 ;
  LAYER metal4 ;
  RECT 1128.460 178.640 1129.580 179.760 ;
  LAYER metal3 ;
  RECT 1128.460 178.640 1129.580 179.760 ;
  LAYER metal2 ;
  RECT 1128.460 178.640 1129.580 179.760 ;
  LAYER metal1 ;
  RECT 1128.460 178.640 1129.580 179.760 ;
 END
END DIB41
PIN DOB41
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1114.820 178.640 1115.940 179.760 ;
  LAYER metal4 ;
  RECT 1114.820 178.640 1115.940 179.760 ;
  LAYER metal3 ;
  RECT 1114.820 178.640 1115.940 179.760 ;
  LAYER metal2 ;
  RECT 1114.820 178.640 1115.940 179.760 ;
  LAYER metal1 ;
  RECT 1114.820 178.640 1115.940 179.760 ;
 END
END DOB41
PIN DIB40
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1101.180 178.640 1102.300 179.760 ;
  LAYER metal4 ;
  RECT 1101.180 178.640 1102.300 179.760 ;
  LAYER metal3 ;
  RECT 1101.180 178.640 1102.300 179.760 ;
  LAYER metal2 ;
  RECT 1101.180 178.640 1102.300 179.760 ;
  LAYER metal1 ;
  RECT 1101.180 178.640 1102.300 179.760 ;
 END
END DIB40
PIN DOB40
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1088.160 178.640 1089.280 179.760 ;
  LAYER metal4 ;
  RECT 1088.160 178.640 1089.280 179.760 ;
  LAYER metal3 ;
  RECT 1088.160 178.640 1089.280 179.760 ;
  LAYER metal2 ;
  RECT 1088.160 178.640 1089.280 179.760 ;
  LAYER metal1 ;
  RECT 1088.160 178.640 1089.280 179.760 ;
 END
END DOB40
PIN DIB39
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1074.520 178.640 1075.640 179.760 ;
  LAYER metal4 ;
  RECT 1074.520 178.640 1075.640 179.760 ;
  LAYER metal3 ;
  RECT 1074.520 178.640 1075.640 179.760 ;
  LAYER metal2 ;
  RECT 1074.520 178.640 1075.640 179.760 ;
  LAYER metal1 ;
  RECT 1074.520 178.640 1075.640 179.760 ;
 END
END DIB39
PIN DOB39
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1060.880 178.640 1062.000 179.760 ;
  LAYER metal4 ;
  RECT 1060.880 178.640 1062.000 179.760 ;
  LAYER metal3 ;
  RECT 1060.880 178.640 1062.000 179.760 ;
  LAYER metal2 ;
  RECT 1060.880 178.640 1062.000 179.760 ;
  LAYER metal1 ;
  RECT 1060.880 178.640 1062.000 179.760 ;
 END
END DOB39
PIN DIB38
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1047.860 178.640 1048.980 179.760 ;
  LAYER metal4 ;
  RECT 1047.860 178.640 1048.980 179.760 ;
  LAYER metal3 ;
  RECT 1047.860 178.640 1048.980 179.760 ;
  LAYER metal2 ;
  RECT 1047.860 178.640 1048.980 179.760 ;
  LAYER metal1 ;
  RECT 1047.860 178.640 1048.980 179.760 ;
 END
END DIB38
PIN DOB38
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1034.220 178.640 1035.340 179.760 ;
  LAYER metal4 ;
  RECT 1034.220 178.640 1035.340 179.760 ;
  LAYER metal3 ;
  RECT 1034.220 178.640 1035.340 179.760 ;
  LAYER metal2 ;
  RECT 1034.220 178.640 1035.340 179.760 ;
  LAYER metal1 ;
  RECT 1034.220 178.640 1035.340 179.760 ;
 END
END DOB38
PIN DIB37
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1020.580 178.640 1021.700 179.760 ;
  LAYER metal4 ;
  RECT 1020.580 178.640 1021.700 179.760 ;
  LAYER metal3 ;
  RECT 1020.580 178.640 1021.700 179.760 ;
  LAYER metal2 ;
  RECT 1020.580 178.640 1021.700 179.760 ;
  LAYER metal1 ;
  RECT 1020.580 178.640 1021.700 179.760 ;
 END
END DIB37
PIN DOB37
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1007.560 178.640 1008.680 179.760 ;
  LAYER metal4 ;
  RECT 1007.560 178.640 1008.680 179.760 ;
  LAYER metal3 ;
  RECT 1007.560 178.640 1008.680 179.760 ;
  LAYER metal2 ;
  RECT 1007.560 178.640 1008.680 179.760 ;
  LAYER metal1 ;
  RECT 1007.560 178.640 1008.680 179.760 ;
 END
END DOB37
PIN DIB36
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 993.920 178.640 995.040 179.760 ;
  LAYER metal4 ;
  RECT 993.920 178.640 995.040 179.760 ;
  LAYER metal3 ;
  RECT 993.920 178.640 995.040 179.760 ;
  LAYER metal2 ;
  RECT 993.920 178.640 995.040 179.760 ;
  LAYER metal1 ;
  RECT 993.920 178.640 995.040 179.760 ;
 END
END DIB36
PIN DOB36
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 980.280 178.640 981.400 179.760 ;
  LAYER metal4 ;
  RECT 980.280 178.640 981.400 179.760 ;
  LAYER metal3 ;
  RECT 980.280 178.640 981.400 179.760 ;
  LAYER metal2 ;
  RECT 980.280 178.640 981.400 179.760 ;
  LAYER metal1 ;
  RECT 980.280 178.640 981.400 179.760 ;
 END
END DOB36
PIN DIB35
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 967.260 178.640 968.380 179.760 ;
  LAYER metal4 ;
  RECT 967.260 178.640 968.380 179.760 ;
  LAYER metal3 ;
  RECT 967.260 178.640 968.380 179.760 ;
  LAYER metal2 ;
  RECT 967.260 178.640 968.380 179.760 ;
  LAYER metal1 ;
  RECT 967.260 178.640 968.380 179.760 ;
 END
END DIB35
PIN DOB35
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 953.620 178.640 954.740 179.760 ;
  LAYER metal4 ;
  RECT 953.620 178.640 954.740 179.760 ;
  LAYER metal3 ;
  RECT 953.620 178.640 954.740 179.760 ;
  LAYER metal2 ;
  RECT 953.620 178.640 954.740 179.760 ;
  LAYER metal1 ;
  RECT 953.620 178.640 954.740 179.760 ;
 END
END DOB35
PIN DIB34
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 939.980 178.640 941.100 179.760 ;
  LAYER metal4 ;
  RECT 939.980 178.640 941.100 179.760 ;
  LAYER metal3 ;
  RECT 939.980 178.640 941.100 179.760 ;
  LAYER metal2 ;
  RECT 939.980 178.640 941.100 179.760 ;
  LAYER metal1 ;
  RECT 939.980 178.640 941.100 179.760 ;
 END
END DIB34
PIN DOB34
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 926.960 178.640 928.080 179.760 ;
  LAYER metal4 ;
  RECT 926.960 178.640 928.080 179.760 ;
  LAYER metal3 ;
  RECT 926.960 178.640 928.080 179.760 ;
  LAYER metal2 ;
  RECT 926.960 178.640 928.080 179.760 ;
  LAYER metal1 ;
  RECT 926.960 178.640 928.080 179.760 ;
 END
END DOB34
PIN DIB33
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 913.320 178.640 914.440 179.760 ;
  LAYER metal4 ;
  RECT 913.320 178.640 914.440 179.760 ;
  LAYER metal3 ;
  RECT 913.320 178.640 914.440 179.760 ;
  LAYER metal2 ;
  RECT 913.320 178.640 914.440 179.760 ;
  LAYER metal1 ;
  RECT 913.320 178.640 914.440 179.760 ;
 END
END DIB33
PIN DOB33
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 899.680 178.640 900.800 179.760 ;
  LAYER metal4 ;
  RECT 899.680 178.640 900.800 179.760 ;
  LAYER metal3 ;
  RECT 899.680 178.640 900.800 179.760 ;
  LAYER metal2 ;
  RECT 899.680 178.640 900.800 179.760 ;
  LAYER metal1 ;
  RECT 899.680 178.640 900.800 179.760 ;
 END
END DOB33
PIN DIB32
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 886.040 178.640 887.160 179.760 ;
  LAYER metal4 ;
  RECT 886.040 178.640 887.160 179.760 ;
  LAYER metal3 ;
  RECT 886.040 178.640 887.160 179.760 ;
  LAYER metal2 ;
  RECT 886.040 178.640 887.160 179.760 ;
  LAYER metal1 ;
  RECT 886.040 178.640 887.160 179.760 ;
 END
END DIB32
PIN WEBN2
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 874.880 178.640 876.000 179.760 ;
  LAYER metal4 ;
  RECT 874.880 178.640 876.000 179.760 ;
  LAYER metal3 ;
  RECT 874.880 178.640 876.000 179.760 ;
  LAYER metal2 ;
  RECT 874.880 178.640 876.000 179.760 ;
  LAYER metal1 ;
  RECT 874.880 178.640 876.000 179.760 ;
 END
END WEBN2
PIN DOB32
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 873.020 178.640 874.140 179.760 ;
  LAYER metal4 ;
  RECT 873.020 178.640 874.140 179.760 ;
  LAYER metal3 ;
  RECT 873.020 178.640 874.140 179.760 ;
  LAYER metal2 ;
  RECT 873.020 178.640 874.140 179.760 ;
  LAYER metal1 ;
  RECT 873.020 178.640 874.140 179.760 ;
 END
END DOB32
PIN DIB31
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 859.380 178.640 860.500 179.760 ;
  LAYER metal4 ;
  RECT 859.380 178.640 860.500 179.760 ;
  LAYER metal3 ;
  RECT 859.380 178.640 860.500 179.760 ;
  LAYER metal2 ;
  RECT 859.380 178.640 860.500 179.760 ;
  LAYER metal1 ;
  RECT 859.380 178.640 860.500 179.760 ;
 END
END DIB31
PIN DOB31
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 845.740 178.640 846.860 179.760 ;
  LAYER metal4 ;
  RECT 845.740 178.640 846.860 179.760 ;
  LAYER metal3 ;
  RECT 845.740 178.640 846.860 179.760 ;
  LAYER metal2 ;
  RECT 845.740 178.640 846.860 179.760 ;
  LAYER metal1 ;
  RECT 845.740 178.640 846.860 179.760 ;
 END
END DOB31
PIN DIB30
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 832.720 178.640 833.840 179.760 ;
  LAYER metal4 ;
  RECT 832.720 178.640 833.840 179.760 ;
  LAYER metal3 ;
  RECT 832.720 178.640 833.840 179.760 ;
  LAYER metal2 ;
  RECT 832.720 178.640 833.840 179.760 ;
  LAYER metal1 ;
  RECT 832.720 178.640 833.840 179.760 ;
 END
END DIB30
PIN DOB30
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 819.080 178.640 820.200 179.760 ;
  LAYER metal4 ;
  RECT 819.080 178.640 820.200 179.760 ;
  LAYER metal3 ;
  RECT 819.080 178.640 820.200 179.760 ;
  LAYER metal2 ;
  RECT 819.080 178.640 820.200 179.760 ;
  LAYER metal1 ;
  RECT 819.080 178.640 820.200 179.760 ;
 END
END DOB30
PIN DIB29
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 805.440 178.640 806.560 179.760 ;
  LAYER metal4 ;
  RECT 805.440 178.640 806.560 179.760 ;
  LAYER metal3 ;
  RECT 805.440 178.640 806.560 179.760 ;
  LAYER metal2 ;
  RECT 805.440 178.640 806.560 179.760 ;
  LAYER metal1 ;
  RECT 805.440 178.640 806.560 179.760 ;
 END
END DIB29
PIN DOB29
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 792.420 178.640 793.540 179.760 ;
  LAYER metal4 ;
  RECT 792.420 178.640 793.540 179.760 ;
  LAYER metal3 ;
  RECT 792.420 178.640 793.540 179.760 ;
  LAYER metal2 ;
  RECT 792.420 178.640 793.540 179.760 ;
  LAYER metal1 ;
  RECT 792.420 178.640 793.540 179.760 ;
 END
END DOB29
PIN DIB28
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 778.780 178.640 779.900 179.760 ;
  LAYER metal4 ;
  RECT 778.780 178.640 779.900 179.760 ;
  LAYER metal3 ;
  RECT 778.780 178.640 779.900 179.760 ;
  LAYER metal2 ;
  RECT 778.780 178.640 779.900 179.760 ;
  LAYER metal1 ;
  RECT 778.780 178.640 779.900 179.760 ;
 END
END DIB28
PIN DOB28
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 765.140 178.640 766.260 179.760 ;
  LAYER metal4 ;
  RECT 765.140 178.640 766.260 179.760 ;
  LAYER metal3 ;
  RECT 765.140 178.640 766.260 179.760 ;
  LAYER metal2 ;
  RECT 765.140 178.640 766.260 179.760 ;
  LAYER metal1 ;
  RECT 765.140 178.640 766.260 179.760 ;
 END
END DOB28
PIN DIB27
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 752.120 178.640 753.240 179.760 ;
  LAYER metal4 ;
  RECT 752.120 178.640 753.240 179.760 ;
  LAYER metal3 ;
  RECT 752.120 178.640 753.240 179.760 ;
  LAYER metal2 ;
  RECT 752.120 178.640 753.240 179.760 ;
  LAYER metal1 ;
  RECT 752.120 178.640 753.240 179.760 ;
 END
END DIB27
PIN DOB27
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 738.480 178.640 739.600 179.760 ;
  LAYER metal4 ;
  RECT 738.480 178.640 739.600 179.760 ;
  LAYER metal3 ;
  RECT 738.480 178.640 739.600 179.760 ;
  LAYER metal2 ;
  RECT 738.480 178.640 739.600 179.760 ;
  LAYER metal1 ;
  RECT 738.480 178.640 739.600 179.760 ;
 END
END DOB27
PIN DIB26
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 724.840 178.640 725.960 179.760 ;
  LAYER metal4 ;
  RECT 724.840 178.640 725.960 179.760 ;
  LAYER metal3 ;
  RECT 724.840 178.640 725.960 179.760 ;
  LAYER metal2 ;
  RECT 724.840 178.640 725.960 179.760 ;
  LAYER metal1 ;
  RECT 724.840 178.640 725.960 179.760 ;
 END
END DIB26
PIN DOB26
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 711.820 178.640 712.940 179.760 ;
  LAYER metal4 ;
  RECT 711.820 178.640 712.940 179.760 ;
  LAYER metal3 ;
  RECT 711.820 178.640 712.940 179.760 ;
  LAYER metal2 ;
  RECT 711.820 178.640 712.940 179.760 ;
  LAYER metal1 ;
  RECT 711.820 178.640 712.940 179.760 ;
 END
END DOB26
PIN DIB25
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 698.180 178.640 699.300 179.760 ;
  LAYER metal4 ;
  RECT 698.180 178.640 699.300 179.760 ;
  LAYER metal3 ;
  RECT 698.180 178.640 699.300 179.760 ;
  LAYER metal2 ;
  RECT 698.180 178.640 699.300 179.760 ;
  LAYER metal1 ;
  RECT 698.180 178.640 699.300 179.760 ;
 END
END DIB25
PIN DOB25
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 684.540 178.640 685.660 179.760 ;
  LAYER metal4 ;
  RECT 684.540 178.640 685.660 179.760 ;
  LAYER metal3 ;
  RECT 684.540 178.640 685.660 179.760 ;
  LAYER metal2 ;
  RECT 684.540 178.640 685.660 179.760 ;
  LAYER metal1 ;
  RECT 684.540 178.640 685.660 179.760 ;
 END
END DOB25
PIN DIB24
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 671.520 178.640 672.640 179.760 ;
  LAYER metal4 ;
  RECT 671.520 178.640 672.640 179.760 ;
  LAYER metal3 ;
  RECT 671.520 178.640 672.640 179.760 ;
  LAYER metal2 ;
  RECT 671.520 178.640 672.640 179.760 ;
  LAYER metal1 ;
  RECT 671.520 178.640 672.640 179.760 ;
 END
END DIB24
PIN DOB24
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 657.880 178.640 659.000 179.760 ;
  LAYER metal4 ;
  RECT 657.880 178.640 659.000 179.760 ;
  LAYER metal3 ;
  RECT 657.880 178.640 659.000 179.760 ;
  LAYER metal2 ;
  RECT 657.880 178.640 659.000 179.760 ;
  LAYER metal1 ;
  RECT 657.880 178.640 659.000 179.760 ;
 END
END DOB24
PIN DIB23
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 644.240 178.640 645.360 179.760 ;
  LAYER metal4 ;
  RECT 644.240 178.640 645.360 179.760 ;
  LAYER metal3 ;
  RECT 644.240 178.640 645.360 179.760 ;
  LAYER metal2 ;
  RECT 644.240 178.640 645.360 179.760 ;
  LAYER metal1 ;
  RECT 644.240 178.640 645.360 179.760 ;
 END
END DIB23
PIN DOB23
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 631.220 178.640 632.340 179.760 ;
  LAYER metal4 ;
  RECT 631.220 178.640 632.340 179.760 ;
  LAYER metal3 ;
  RECT 631.220 178.640 632.340 179.760 ;
  LAYER metal2 ;
  RECT 631.220 178.640 632.340 179.760 ;
  LAYER metal1 ;
  RECT 631.220 178.640 632.340 179.760 ;
 END
END DOB23
PIN DIB22
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 617.580 178.640 618.700 179.760 ;
  LAYER metal4 ;
  RECT 617.580 178.640 618.700 179.760 ;
  LAYER metal3 ;
  RECT 617.580 178.640 618.700 179.760 ;
  LAYER metal2 ;
  RECT 617.580 178.640 618.700 179.760 ;
  LAYER metal1 ;
  RECT 617.580 178.640 618.700 179.760 ;
 END
END DIB22
PIN DOB22
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 603.940 178.640 605.060 179.760 ;
  LAYER metal4 ;
  RECT 603.940 178.640 605.060 179.760 ;
  LAYER metal3 ;
  RECT 603.940 178.640 605.060 179.760 ;
  LAYER metal2 ;
  RECT 603.940 178.640 605.060 179.760 ;
  LAYER metal1 ;
  RECT 603.940 178.640 605.060 179.760 ;
 END
END DOB22
PIN DIB21
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 590.920 178.640 592.040 179.760 ;
  LAYER metal4 ;
  RECT 590.920 178.640 592.040 179.760 ;
  LAYER metal3 ;
  RECT 590.920 178.640 592.040 179.760 ;
  LAYER metal2 ;
  RECT 590.920 178.640 592.040 179.760 ;
  LAYER metal1 ;
  RECT 590.920 178.640 592.040 179.760 ;
 END
END DIB21
PIN DOB21
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 577.280 178.640 578.400 179.760 ;
  LAYER metal4 ;
  RECT 577.280 178.640 578.400 179.760 ;
  LAYER metal3 ;
  RECT 577.280 178.640 578.400 179.760 ;
  LAYER metal2 ;
  RECT 577.280 178.640 578.400 179.760 ;
  LAYER metal1 ;
  RECT 577.280 178.640 578.400 179.760 ;
 END
END DOB21
PIN DIB20
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 563.640 178.640 564.760 179.760 ;
  LAYER metal4 ;
  RECT 563.640 178.640 564.760 179.760 ;
  LAYER metal3 ;
  RECT 563.640 178.640 564.760 179.760 ;
  LAYER metal2 ;
  RECT 563.640 178.640 564.760 179.760 ;
  LAYER metal1 ;
  RECT 563.640 178.640 564.760 179.760 ;
 END
END DIB20
PIN DOB20
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 550.620 178.640 551.740 179.760 ;
  LAYER metal4 ;
  RECT 550.620 178.640 551.740 179.760 ;
  LAYER metal3 ;
  RECT 550.620 178.640 551.740 179.760 ;
  LAYER metal2 ;
  RECT 550.620 178.640 551.740 179.760 ;
  LAYER metal1 ;
  RECT 550.620 178.640 551.740 179.760 ;
 END
END DOB20
PIN DIB19
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 536.980 178.640 538.100 179.760 ;
  LAYER metal4 ;
  RECT 536.980 178.640 538.100 179.760 ;
  LAYER metal3 ;
  RECT 536.980 178.640 538.100 179.760 ;
  LAYER metal2 ;
  RECT 536.980 178.640 538.100 179.760 ;
  LAYER metal1 ;
  RECT 536.980 178.640 538.100 179.760 ;
 END
END DIB19
PIN DOB19
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 523.340 178.640 524.460 179.760 ;
  LAYER metal4 ;
  RECT 523.340 178.640 524.460 179.760 ;
  LAYER metal3 ;
  RECT 523.340 178.640 524.460 179.760 ;
  LAYER metal2 ;
  RECT 523.340 178.640 524.460 179.760 ;
  LAYER metal1 ;
  RECT 523.340 178.640 524.460 179.760 ;
 END
END DOB19
PIN DIB18
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 510.320 178.640 511.440 179.760 ;
  LAYER metal4 ;
  RECT 510.320 178.640 511.440 179.760 ;
  LAYER metal3 ;
  RECT 510.320 178.640 511.440 179.760 ;
  LAYER metal2 ;
  RECT 510.320 178.640 511.440 179.760 ;
  LAYER metal1 ;
  RECT 510.320 178.640 511.440 179.760 ;
 END
END DIB18
PIN DOB18
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 496.680 178.640 497.800 179.760 ;
  LAYER metal4 ;
  RECT 496.680 178.640 497.800 179.760 ;
  LAYER metal3 ;
  RECT 496.680 178.640 497.800 179.760 ;
  LAYER metal2 ;
  RECT 496.680 178.640 497.800 179.760 ;
  LAYER metal1 ;
  RECT 496.680 178.640 497.800 179.760 ;
 END
END DOB18
PIN DIB17
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 483.040 178.640 484.160 179.760 ;
  LAYER metal4 ;
  RECT 483.040 178.640 484.160 179.760 ;
  LAYER metal3 ;
  RECT 483.040 178.640 484.160 179.760 ;
  LAYER metal2 ;
  RECT 483.040 178.640 484.160 179.760 ;
  LAYER metal1 ;
  RECT 483.040 178.640 484.160 179.760 ;
 END
END DIB17
PIN DOB17
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 469.400 178.640 470.520 179.760 ;
  LAYER metal4 ;
  RECT 469.400 178.640 470.520 179.760 ;
  LAYER metal3 ;
  RECT 469.400 178.640 470.520 179.760 ;
  LAYER metal2 ;
  RECT 469.400 178.640 470.520 179.760 ;
  LAYER metal1 ;
  RECT 469.400 178.640 470.520 179.760 ;
 END
END DOB17
PIN DIB16
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 456.380 178.640 457.500 179.760 ;
  LAYER metal4 ;
  RECT 456.380 178.640 457.500 179.760 ;
  LAYER metal3 ;
  RECT 456.380 178.640 457.500 179.760 ;
  LAYER metal2 ;
  RECT 456.380 178.640 457.500 179.760 ;
  LAYER metal1 ;
  RECT 456.380 178.640 457.500 179.760 ;
 END
END DIB16
PIN WEBN1
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 445.220 178.640 446.340 179.760 ;
  LAYER metal4 ;
  RECT 445.220 178.640 446.340 179.760 ;
  LAYER metal3 ;
  RECT 445.220 178.640 446.340 179.760 ;
  LAYER metal2 ;
  RECT 445.220 178.640 446.340 179.760 ;
  LAYER metal1 ;
  RECT 445.220 178.640 446.340 179.760 ;
 END
END WEBN1
PIN DOB16
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 442.740 178.640 443.860 179.760 ;
  LAYER metal4 ;
  RECT 442.740 178.640 443.860 179.760 ;
  LAYER metal3 ;
  RECT 442.740 178.640 443.860 179.760 ;
  LAYER metal2 ;
  RECT 442.740 178.640 443.860 179.760 ;
  LAYER metal1 ;
  RECT 442.740 178.640 443.860 179.760 ;
 END
END DOB16
PIN DIB15
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 429.100 178.640 430.220 179.760 ;
  LAYER metal4 ;
  RECT 429.100 178.640 430.220 179.760 ;
  LAYER metal3 ;
  RECT 429.100 178.640 430.220 179.760 ;
  LAYER metal2 ;
  RECT 429.100 178.640 430.220 179.760 ;
  LAYER metal1 ;
  RECT 429.100 178.640 430.220 179.760 ;
 END
END DIB15
PIN DOB15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 416.080 178.640 417.200 179.760 ;
  LAYER metal4 ;
  RECT 416.080 178.640 417.200 179.760 ;
  LAYER metal3 ;
  RECT 416.080 178.640 417.200 179.760 ;
  LAYER metal2 ;
  RECT 416.080 178.640 417.200 179.760 ;
  LAYER metal1 ;
  RECT 416.080 178.640 417.200 179.760 ;
 END
END DOB15
PIN DIB14
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 402.440 178.640 403.560 179.760 ;
  LAYER metal4 ;
  RECT 402.440 178.640 403.560 179.760 ;
  LAYER metal3 ;
  RECT 402.440 178.640 403.560 179.760 ;
  LAYER metal2 ;
  RECT 402.440 178.640 403.560 179.760 ;
  LAYER metal1 ;
  RECT 402.440 178.640 403.560 179.760 ;
 END
END DIB14
PIN DOB14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 388.800 178.640 389.920 179.760 ;
  LAYER metal4 ;
  RECT 388.800 178.640 389.920 179.760 ;
  LAYER metal3 ;
  RECT 388.800 178.640 389.920 179.760 ;
  LAYER metal2 ;
  RECT 388.800 178.640 389.920 179.760 ;
  LAYER metal1 ;
  RECT 388.800 178.640 389.920 179.760 ;
 END
END DOB14
PIN DIB13
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 375.780 178.640 376.900 179.760 ;
  LAYER metal4 ;
  RECT 375.780 178.640 376.900 179.760 ;
  LAYER metal3 ;
  RECT 375.780 178.640 376.900 179.760 ;
  LAYER metal2 ;
  RECT 375.780 178.640 376.900 179.760 ;
  LAYER metal1 ;
  RECT 375.780 178.640 376.900 179.760 ;
 END
END DIB13
PIN DOB13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 362.140 178.640 363.260 179.760 ;
  LAYER metal4 ;
  RECT 362.140 178.640 363.260 179.760 ;
  LAYER metal3 ;
  RECT 362.140 178.640 363.260 179.760 ;
  LAYER metal2 ;
  RECT 362.140 178.640 363.260 179.760 ;
  LAYER metal1 ;
  RECT 362.140 178.640 363.260 179.760 ;
 END
END DOB13
PIN DIB12
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 348.500 178.640 349.620 179.760 ;
  LAYER metal4 ;
  RECT 348.500 178.640 349.620 179.760 ;
  LAYER metal3 ;
  RECT 348.500 178.640 349.620 179.760 ;
  LAYER metal2 ;
  RECT 348.500 178.640 349.620 179.760 ;
  LAYER metal1 ;
  RECT 348.500 178.640 349.620 179.760 ;
 END
END DIB12
PIN DOB12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 335.480 178.640 336.600 179.760 ;
  LAYER metal4 ;
  RECT 335.480 178.640 336.600 179.760 ;
  LAYER metal3 ;
  RECT 335.480 178.640 336.600 179.760 ;
  LAYER metal2 ;
  RECT 335.480 178.640 336.600 179.760 ;
  LAYER metal1 ;
  RECT 335.480 178.640 336.600 179.760 ;
 END
END DOB12
PIN DIB11
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 321.840 178.640 322.960 179.760 ;
  LAYER metal4 ;
  RECT 321.840 178.640 322.960 179.760 ;
  LAYER metal3 ;
  RECT 321.840 178.640 322.960 179.760 ;
  LAYER metal2 ;
  RECT 321.840 178.640 322.960 179.760 ;
  LAYER metal1 ;
  RECT 321.840 178.640 322.960 179.760 ;
 END
END DIB11
PIN DOB11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 308.200 178.640 309.320 179.760 ;
  LAYER metal4 ;
  RECT 308.200 178.640 309.320 179.760 ;
  LAYER metal3 ;
  RECT 308.200 178.640 309.320 179.760 ;
  LAYER metal2 ;
  RECT 308.200 178.640 309.320 179.760 ;
  LAYER metal1 ;
  RECT 308.200 178.640 309.320 179.760 ;
 END
END DOB11
PIN DIB10
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 295.180 178.640 296.300 179.760 ;
  LAYER metal4 ;
  RECT 295.180 178.640 296.300 179.760 ;
  LAYER metal3 ;
  RECT 295.180 178.640 296.300 179.760 ;
  LAYER metal2 ;
  RECT 295.180 178.640 296.300 179.760 ;
  LAYER metal1 ;
  RECT 295.180 178.640 296.300 179.760 ;
 END
END DIB10
PIN DOB10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 281.540 178.640 282.660 179.760 ;
  LAYER metal4 ;
  RECT 281.540 178.640 282.660 179.760 ;
  LAYER metal3 ;
  RECT 281.540 178.640 282.660 179.760 ;
  LAYER metal2 ;
  RECT 281.540 178.640 282.660 179.760 ;
  LAYER metal1 ;
  RECT 281.540 178.640 282.660 179.760 ;
 END
END DOB10
PIN DIB9
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 267.900 178.640 269.020 179.760 ;
  LAYER metal4 ;
  RECT 267.900 178.640 269.020 179.760 ;
  LAYER metal3 ;
  RECT 267.900 178.640 269.020 179.760 ;
  LAYER metal2 ;
  RECT 267.900 178.640 269.020 179.760 ;
  LAYER metal1 ;
  RECT 267.900 178.640 269.020 179.760 ;
 END
END DIB9
PIN DOB9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 254.880 178.640 256.000 179.760 ;
  LAYER metal4 ;
  RECT 254.880 178.640 256.000 179.760 ;
  LAYER metal3 ;
  RECT 254.880 178.640 256.000 179.760 ;
  LAYER metal2 ;
  RECT 254.880 178.640 256.000 179.760 ;
  LAYER metal1 ;
  RECT 254.880 178.640 256.000 179.760 ;
 END
END DOB9
PIN DIB8
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 241.240 178.640 242.360 179.760 ;
  LAYER metal4 ;
  RECT 241.240 178.640 242.360 179.760 ;
  LAYER metal3 ;
  RECT 241.240 178.640 242.360 179.760 ;
  LAYER metal2 ;
  RECT 241.240 178.640 242.360 179.760 ;
  LAYER metal1 ;
  RECT 241.240 178.640 242.360 179.760 ;
 END
END DIB8
PIN DOB8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 227.600 178.640 228.720 179.760 ;
  LAYER metal4 ;
  RECT 227.600 178.640 228.720 179.760 ;
  LAYER metal3 ;
  RECT 227.600 178.640 228.720 179.760 ;
  LAYER metal2 ;
  RECT 227.600 178.640 228.720 179.760 ;
  LAYER metal1 ;
  RECT 227.600 178.640 228.720 179.760 ;
 END
END DOB8
PIN DIB7
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 214.580 178.640 215.700 179.760 ;
  LAYER metal4 ;
  RECT 214.580 178.640 215.700 179.760 ;
  LAYER metal3 ;
  RECT 214.580 178.640 215.700 179.760 ;
  LAYER metal2 ;
  RECT 214.580 178.640 215.700 179.760 ;
  LAYER metal1 ;
  RECT 214.580 178.640 215.700 179.760 ;
 END
END DIB7
PIN DOB7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 200.940 178.640 202.060 179.760 ;
  LAYER metal4 ;
  RECT 200.940 178.640 202.060 179.760 ;
  LAYER metal3 ;
  RECT 200.940 178.640 202.060 179.760 ;
  LAYER metal2 ;
  RECT 200.940 178.640 202.060 179.760 ;
  LAYER metal1 ;
  RECT 200.940 178.640 202.060 179.760 ;
 END
END DOB7
PIN DIB6
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 187.300 178.640 188.420 179.760 ;
  LAYER metal4 ;
  RECT 187.300 178.640 188.420 179.760 ;
  LAYER metal3 ;
  RECT 187.300 178.640 188.420 179.760 ;
  LAYER metal2 ;
  RECT 187.300 178.640 188.420 179.760 ;
  LAYER metal1 ;
  RECT 187.300 178.640 188.420 179.760 ;
 END
END DIB6
PIN DOB6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 174.280 178.640 175.400 179.760 ;
  LAYER metal4 ;
  RECT 174.280 178.640 175.400 179.760 ;
  LAYER metal3 ;
  RECT 174.280 178.640 175.400 179.760 ;
  LAYER metal2 ;
  RECT 174.280 178.640 175.400 179.760 ;
  LAYER metal1 ;
  RECT 174.280 178.640 175.400 179.760 ;
 END
END DOB6
PIN DIB5
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 160.640 178.640 161.760 179.760 ;
  LAYER metal4 ;
  RECT 160.640 178.640 161.760 179.760 ;
  LAYER metal3 ;
  RECT 160.640 178.640 161.760 179.760 ;
  LAYER metal2 ;
  RECT 160.640 178.640 161.760 179.760 ;
  LAYER metal1 ;
  RECT 160.640 178.640 161.760 179.760 ;
 END
END DIB5
PIN DOB5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 147.000 178.640 148.120 179.760 ;
  LAYER metal4 ;
  RECT 147.000 178.640 148.120 179.760 ;
  LAYER metal3 ;
  RECT 147.000 178.640 148.120 179.760 ;
  LAYER metal2 ;
  RECT 147.000 178.640 148.120 179.760 ;
  LAYER metal1 ;
  RECT 147.000 178.640 148.120 179.760 ;
 END
END DOB5
PIN DIB4
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 133.980 178.640 135.100 179.760 ;
  LAYER metal4 ;
  RECT 133.980 178.640 135.100 179.760 ;
  LAYER metal3 ;
  RECT 133.980 178.640 135.100 179.760 ;
  LAYER metal2 ;
  RECT 133.980 178.640 135.100 179.760 ;
  LAYER metal1 ;
  RECT 133.980 178.640 135.100 179.760 ;
 END
END DIB4
PIN DOB4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 120.340 178.640 121.460 179.760 ;
  LAYER metal4 ;
  RECT 120.340 178.640 121.460 179.760 ;
  LAYER metal3 ;
  RECT 120.340 178.640 121.460 179.760 ;
  LAYER metal2 ;
  RECT 120.340 178.640 121.460 179.760 ;
  LAYER metal1 ;
  RECT 120.340 178.640 121.460 179.760 ;
 END
END DOB4
PIN DIB3
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 106.700 178.640 107.820 179.760 ;
  LAYER metal4 ;
  RECT 106.700 178.640 107.820 179.760 ;
  LAYER metal3 ;
  RECT 106.700 178.640 107.820 179.760 ;
  LAYER metal2 ;
  RECT 106.700 178.640 107.820 179.760 ;
  LAYER metal1 ;
  RECT 106.700 178.640 107.820 179.760 ;
 END
END DIB3
PIN DOB3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 93.680 178.640 94.800 179.760 ;
  LAYER metal4 ;
  RECT 93.680 178.640 94.800 179.760 ;
  LAYER metal3 ;
  RECT 93.680 178.640 94.800 179.760 ;
  LAYER metal2 ;
  RECT 93.680 178.640 94.800 179.760 ;
  LAYER metal1 ;
  RECT 93.680 178.640 94.800 179.760 ;
 END
END DOB3
PIN DIB2
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 80.040 178.640 81.160 179.760 ;
  LAYER metal4 ;
  RECT 80.040 178.640 81.160 179.760 ;
  LAYER metal3 ;
  RECT 80.040 178.640 81.160 179.760 ;
  LAYER metal2 ;
  RECT 80.040 178.640 81.160 179.760 ;
  LAYER metal1 ;
  RECT 80.040 178.640 81.160 179.760 ;
 END
END DIB2
PIN DOB2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 66.400 178.640 67.520 179.760 ;
  LAYER metal4 ;
  RECT 66.400 178.640 67.520 179.760 ;
  LAYER metal3 ;
  RECT 66.400 178.640 67.520 179.760 ;
  LAYER metal2 ;
  RECT 66.400 178.640 67.520 179.760 ;
  LAYER metal1 ;
  RECT 66.400 178.640 67.520 179.760 ;
 END
END DOB2
PIN DIB1
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 52.760 178.640 53.880 179.760 ;
  LAYER metal4 ;
  RECT 52.760 178.640 53.880 179.760 ;
  LAYER metal3 ;
  RECT 52.760 178.640 53.880 179.760 ;
  LAYER metal2 ;
  RECT 52.760 178.640 53.880 179.760 ;
  LAYER metal1 ;
  RECT 52.760 178.640 53.880 179.760 ;
 END
END DIB1
PIN DOB1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 39.740 178.640 40.860 179.760 ;
  LAYER metal4 ;
  RECT 39.740 178.640 40.860 179.760 ;
  LAYER metal3 ;
  RECT 39.740 178.640 40.860 179.760 ;
  LAYER metal2 ;
  RECT 39.740 178.640 40.860 179.760 ;
  LAYER metal1 ;
  RECT 39.740 178.640 40.860 179.760 ;
 END
END DOB1
PIN DIB0
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 26.100 178.640 27.220 179.760 ;
  LAYER metal4 ;
  RECT 26.100 178.640 27.220 179.760 ;
  LAYER metal3 ;
  RECT 26.100 178.640 27.220 179.760 ;
  LAYER metal2 ;
  RECT 26.100 178.640 27.220 179.760 ;
  LAYER metal1 ;
  RECT 26.100 178.640 27.220 179.760 ;
 END
END DIB0
PIN WEBN0
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 14.940 178.640 16.060 179.760 ;
  LAYER metal4 ;
  RECT 14.940 178.640 16.060 179.760 ;
  LAYER metal3 ;
  RECT 14.940 178.640 16.060 179.760 ;
  LAYER metal2 ;
  RECT 14.940 178.640 16.060 179.760 ;
  LAYER metal1 ;
  RECT 14.940 178.640 16.060 179.760 ;
 END
END WEBN0
PIN DOB0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 12.460 178.640 13.580 179.760 ;
  LAYER metal4 ;
  RECT 12.460 178.640 13.580 179.760 ;
  LAYER metal3 ;
  RECT 12.460 178.640 13.580 179.760 ;
  LAYER metal2 ;
  RECT 12.460 178.640 13.580 179.760 ;
  LAYER metal1 ;
  RECT 12.460 178.640 13.580 179.760 ;
 END
END DOB0
PIN DIA127
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3524.760 0.000 3525.880 1.120 ;
  LAYER metal4 ;
  RECT 3524.760 0.000 3525.880 1.120 ;
  LAYER metal3 ;
  RECT 3524.760 0.000 3525.880 1.120 ;
  LAYER metal2 ;
  RECT 3524.760 0.000 3525.880 1.120 ;
  LAYER metal1 ;
  RECT 3524.760 0.000 3525.880 1.120 ;
 END
END DIA127
PIN DOA127
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3511.120 0.000 3512.240 1.120 ;
  LAYER metal4 ;
  RECT 3511.120 0.000 3512.240 1.120 ;
  LAYER metal3 ;
  RECT 3511.120 0.000 3512.240 1.120 ;
  LAYER metal2 ;
  RECT 3511.120 0.000 3512.240 1.120 ;
  LAYER metal1 ;
  RECT 3511.120 0.000 3512.240 1.120 ;
 END
END DOA127
PIN DIA126
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3497.480 0.000 3498.600 1.120 ;
  LAYER metal4 ;
  RECT 3497.480 0.000 3498.600 1.120 ;
  LAYER metal3 ;
  RECT 3497.480 0.000 3498.600 1.120 ;
  LAYER metal2 ;
  RECT 3497.480 0.000 3498.600 1.120 ;
  LAYER metal1 ;
  RECT 3497.480 0.000 3498.600 1.120 ;
 END
END DIA126
PIN DOA126
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3484.460 0.000 3485.580 1.120 ;
  LAYER metal4 ;
  RECT 3484.460 0.000 3485.580 1.120 ;
  LAYER metal3 ;
  RECT 3484.460 0.000 3485.580 1.120 ;
  LAYER metal2 ;
  RECT 3484.460 0.000 3485.580 1.120 ;
  LAYER metal1 ;
  RECT 3484.460 0.000 3485.580 1.120 ;
 END
END DOA126
PIN DIA125
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3470.820 0.000 3471.940 1.120 ;
  LAYER metal4 ;
  RECT 3470.820 0.000 3471.940 1.120 ;
  LAYER metal3 ;
  RECT 3470.820 0.000 3471.940 1.120 ;
  LAYER metal2 ;
  RECT 3470.820 0.000 3471.940 1.120 ;
  LAYER metal1 ;
  RECT 3470.820 0.000 3471.940 1.120 ;
 END
END DIA125
PIN DOA125
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3457.180 0.000 3458.300 1.120 ;
  LAYER metal4 ;
  RECT 3457.180 0.000 3458.300 1.120 ;
  LAYER metal3 ;
  RECT 3457.180 0.000 3458.300 1.120 ;
  LAYER metal2 ;
  RECT 3457.180 0.000 3458.300 1.120 ;
  LAYER metal1 ;
  RECT 3457.180 0.000 3458.300 1.120 ;
 END
END DOA125
PIN DIA124
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3444.160 0.000 3445.280 1.120 ;
  LAYER metal4 ;
  RECT 3444.160 0.000 3445.280 1.120 ;
  LAYER metal3 ;
  RECT 3444.160 0.000 3445.280 1.120 ;
  LAYER metal2 ;
  RECT 3444.160 0.000 3445.280 1.120 ;
  LAYER metal1 ;
  RECT 3444.160 0.000 3445.280 1.120 ;
 END
END DIA124
PIN DOA124
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3430.520 0.000 3431.640 1.120 ;
  LAYER metal4 ;
  RECT 3430.520 0.000 3431.640 1.120 ;
  LAYER metal3 ;
  RECT 3430.520 0.000 3431.640 1.120 ;
  LAYER metal2 ;
  RECT 3430.520 0.000 3431.640 1.120 ;
  LAYER metal1 ;
  RECT 3430.520 0.000 3431.640 1.120 ;
 END
END DOA124
PIN DIA123
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3416.880 0.000 3418.000 1.120 ;
  LAYER metal4 ;
  RECT 3416.880 0.000 3418.000 1.120 ;
  LAYER metal3 ;
  RECT 3416.880 0.000 3418.000 1.120 ;
  LAYER metal2 ;
  RECT 3416.880 0.000 3418.000 1.120 ;
  LAYER metal1 ;
  RECT 3416.880 0.000 3418.000 1.120 ;
 END
END DIA123
PIN DOA123
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3403.860 0.000 3404.980 1.120 ;
  LAYER metal4 ;
  RECT 3403.860 0.000 3404.980 1.120 ;
  LAYER metal3 ;
  RECT 3403.860 0.000 3404.980 1.120 ;
  LAYER metal2 ;
  RECT 3403.860 0.000 3404.980 1.120 ;
  LAYER metal1 ;
  RECT 3403.860 0.000 3404.980 1.120 ;
 END
END DOA123
PIN DIA122
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3390.220 0.000 3391.340 1.120 ;
  LAYER metal4 ;
  RECT 3390.220 0.000 3391.340 1.120 ;
  LAYER metal3 ;
  RECT 3390.220 0.000 3391.340 1.120 ;
  LAYER metal2 ;
  RECT 3390.220 0.000 3391.340 1.120 ;
  LAYER metal1 ;
  RECT 3390.220 0.000 3391.340 1.120 ;
 END
END DIA122
PIN DOA122
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3376.580 0.000 3377.700 1.120 ;
  LAYER metal4 ;
  RECT 3376.580 0.000 3377.700 1.120 ;
  LAYER metal3 ;
  RECT 3376.580 0.000 3377.700 1.120 ;
  LAYER metal2 ;
  RECT 3376.580 0.000 3377.700 1.120 ;
  LAYER metal1 ;
  RECT 3376.580 0.000 3377.700 1.120 ;
 END
END DOA122
PIN DIA121
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3363.560 0.000 3364.680 1.120 ;
  LAYER metal4 ;
  RECT 3363.560 0.000 3364.680 1.120 ;
  LAYER metal3 ;
  RECT 3363.560 0.000 3364.680 1.120 ;
  LAYER metal2 ;
  RECT 3363.560 0.000 3364.680 1.120 ;
  LAYER metal1 ;
  RECT 3363.560 0.000 3364.680 1.120 ;
 END
END DIA121
PIN DOA121
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3349.920 0.000 3351.040 1.120 ;
  LAYER metal4 ;
  RECT 3349.920 0.000 3351.040 1.120 ;
  LAYER metal3 ;
  RECT 3349.920 0.000 3351.040 1.120 ;
  LAYER metal2 ;
  RECT 3349.920 0.000 3351.040 1.120 ;
  LAYER metal1 ;
  RECT 3349.920 0.000 3351.040 1.120 ;
 END
END DOA121
PIN DIA120
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3336.280 0.000 3337.400 1.120 ;
  LAYER metal4 ;
  RECT 3336.280 0.000 3337.400 1.120 ;
  LAYER metal3 ;
  RECT 3336.280 0.000 3337.400 1.120 ;
  LAYER metal2 ;
  RECT 3336.280 0.000 3337.400 1.120 ;
  LAYER metal1 ;
  RECT 3336.280 0.000 3337.400 1.120 ;
 END
END DIA120
PIN DOA120
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3322.640 0.000 3323.760 1.120 ;
  LAYER metal4 ;
  RECT 3322.640 0.000 3323.760 1.120 ;
  LAYER metal3 ;
  RECT 3322.640 0.000 3323.760 1.120 ;
  LAYER metal2 ;
  RECT 3322.640 0.000 3323.760 1.120 ;
  LAYER metal1 ;
  RECT 3322.640 0.000 3323.760 1.120 ;
 END
END DOA120
PIN DIA119
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3309.620 0.000 3310.740 1.120 ;
  LAYER metal4 ;
  RECT 3309.620 0.000 3310.740 1.120 ;
  LAYER metal3 ;
  RECT 3309.620 0.000 3310.740 1.120 ;
  LAYER metal2 ;
  RECT 3309.620 0.000 3310.740 1.120 ;
  LAYER metal1 ;
  RECT 3309.620 0.000 3310.740 1.120 ;
 END
END DIA119
PIN DOA119
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3295.980 0.000 3297.100 1.120 ;
  LAYER metal4 ;
  RECT 3295.980 0.000 3297.100 1.120 ;
  LAYER metal3 ;
  RECT 3295.980 0.000 3297.100 1.120 ;
  LAYER metal2 ;
  RECT 3295.980 0.000 3297.100 1.120 ;
  LAYER metal1 ;
  RECT 3295.980 0.000 3297.100 1.120 ;
 END
END DOA119
PIN DIA118
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3282.340 0.000 3283.460 1.120 ;
  LAYER metal4 ;
  RECT 3282.340 0.000 3283.460 1.120 ;
  LAYER metal3 ;
  RECT 3282.340 0.000 3283.460 1.120 ;
  LAYER metal2 ;
  RECT 3282.340 0.000 3283.460 1.120 ;
  LAYER metal1 ;
  RECT 3282.340 0.000 3283.460 1.120 ;
 END
END DIA118
PIN DOA118
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3269.320 0.000 3270.440 1.120 ;
  LAYER metal4 ;
  RECT 3269.320 0.000 3270.440 1.120 ;
  LAYER metal3 ;
  RECT 3269.320 0.000 3270.440 1.120 ;
  LAYER metal2 ;
  RECT 3269.320 0.000 3270.440 1.120 ;
  LAYER metal1 ;
  RECT 3269.320 0.000 3270.440 1.120 ;
 END
END DOA118
PIN DIA117
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3255.680 0.000 3256.800 1.120 ;
  LAYER metal4 ;
  RECT 3255.680 0.000 3256.800 1.120 ;
  LAYER metal3 ;
  RECT 3255.680 0.000 3256.800 1.120 ;
  LAYER metal2 ;
  RECT 3255.680 0.000 3256.800 1.120 ;
  LAYER metal1 ;
  RECT 3255.680 0.000 3256.800 1.120 ;
 END
END DIA117
PIN DOA117
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3242.040 0.000 3243.160 1.120 ;
  LAYER metal4 ;
  RECT 3242.040 0.000 3243.160 1.120 ;
  LAYER metal3 ;
  RECT 3242.040 0.000 3243.160 1.120 ;
  LAYER metal2 ;
  RECT 3242.040 0.000 3243.160 1.120 ;
  LAYER metal1 ;
  RECT 3242.040 0.000 3243.160 1.120 ;
 END
END DOA117
PIN DIA116
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3229.020 0.000 3230.140 1.120 ;
  LAYER metal4 ;
  RECT 3229.020 0.000 3230.140 1.120 ;
  LAYER metal3 ;
  RECT 3229.020 0.000 3230.140 1.120 ;
  LAYER metal2 ;
  RECT 3229.020 0.000 3230.140 1.120 ;
  LAYER metal1 ;
  RECT 3229.020 0.000 3230.140 1.120 ;
 END
END DIA116
PIN DOA116
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3215.380 0.000 3216.500 1.120 ;
  LAYER metal4 ;
  RECT 3215.380 0.000 3216.500 1.120 ;
  LAYER metal3 ;
  RECT 3215.380 0.000 3216.500 1.120 ;
  LAYER metal2 ;
  RECT 3215.380 0.000 3216.500 1.120 ;
  LAYER metal1 ;
  RECT 3215.380 0.000 3216.500 1.120 ;
 END
END DOA116
PIN DIA115
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3201.740 0.000 3202.860 1.120 ;
  LAYER metal4 ;
  RECT 3201.740 0.000 3202.860 1.120 ;
  LAYER metal3 ;
  RECT 3201.740 0.000 3202.860 1.120 ;
  LAYER metal2 ;
  RECT 3201.740 0.000 3202.860 1.120 ;
  LAYER metal1 ;
  RECT 3201.740 0.000 3202.860 1.120 ;
 END
END DIA115
PIN DOA115
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3188.720 0.000 3189.840 1.120 ;
  LAYER metal4 ;
  RECT 3188.720 0.000 3189.840 1.120 ;
  LAYER metal3 ;
  RECT 3188.720 0.000 3189.840 1.120 ;
  LAYER metal2 ;
  RECT 3188.720 0.000 3189.840 1.120 ;
  LAYER metal1 ;
  RECT 3188.720 0.000 3189.840 1.120 ;
 END
END DOA115
PIN DIA114
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3175.080 0.000 3176.200 1.120 ;
  LAYER metal4 ;
  RECT 3175.080 0.000 3176.200 1.120 ;
  LAYER metal3 ;
  RECT 3175.080 0.000 3176.200 1.120 ;
  LAYER metal2 ;
  RECT 3175.080 0.000 3176.200 1.120 ;
  LAYER metal1 ;
  RECT 3175.080 0.000 3176.200 1.120 ;
 END
END DIA114
PIN DOA114
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3161.440 0.000 3162.560 1.120 ;
  LAYER metal4 ;
  RECT 3161.440 0.000 3162.560 1.120 ;
  LAYER metal3 ;
  RECT 3161.440 0.000 3162.560 1.120 ;
  LAYER metal2 ;
  RECT 3161.440 0.000 3162.560 1.120 ;
  LAYER metal1 ;
  RECT 3161.440 0.000 3162.560 1.120 ;
 END
END DOA114
PIN DIA113
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3148.420 0.000 3149.540 1.120 ;
  LAYER metal4 ;
  RECT 3148.420 0.000 3149.540 1.120 ;
  LAYER metal3 ;
  RECT 3148.420 0.000 3149.540 1.120 ;
  LAYER metal2 ;
  RECT 3148.420 0.000 3149.540 1.120 ;
  LAYER metal1 ;
  RECT 3148.420 0.000 3149.540 1.120 ;
 END
END DIA113
PIN DOA113
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3134.780 0.000 3135.900 1.120 ;
  LAYER metal4 ;
  RECT 3134.780 0.000 3135.900 1.120 ;
  LAYER metal3 ;
  RECT 3134.780 0.000 3135.900 1.120 ;
  LAYER metal2 ;
  RECT 3134.780 0.000 3135.900 1.120 ;
  LAYER metal1 ;
  RECT 3134.780 0.000 3135.900 1.120 ;
 END
END DOA113
PIN DIA112
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3121.140 0.000 3122.260 1.120 ;
  LAYER metal4 ;
  RECT 3121.140 0.000 3122.260 1.120 ;
  LAYER metal3 ;
  RECT 3121.140 0.000 3122.260 1.120 ;
  LAYER metal2 ;
  RECT 3121.140 0.000 3122.260 1.120 ;
  LAYER metal1 ;
  RECT 3121.140 0.000 3122.260 1.120 ;
 END
END DIA112
PIN WEAN7
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 3109.980 0.000 3111.100 1.120 ;
  LAYER metal4 ;
  RECT 3109.980 0.000 3111.100 1.120 ;
  LAYER metal3 ;
  RECT 3109.980 0.000 3111.100 1.120 ;
  LAYER metal2 ;
  RECT 3109.980 0.000 3111.100 1.120 ;
  LAYER metal1 ;
  RECT 3109.980 0.000 3111.100 1.120 ;
 END
END WEAN7
PIN DOA112
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3108.120 0.000 3109.240 1.120 ;
  LAYER metal4 ;
  RECT 3108.120 0.000 3109.240 1.120 ;
  LAYER metal3 ;
  RECT 3108.120 0.000 3109.240 1.120 ;
  LAYER metal2 ;
  RECT 3108.120 0.000 3109.240 1.120 ;
  LAYER metal1 ;
  RECT 3108.120 0.000 3109.240 1.120 ;
 END
END DOA112
PIN DIA111
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3094.480 0.000 3095.600 1.120 ;
  LAYER metal4 ;
  RECT 3094.480 0.000 3095.600 1.120 ;
  LAYER metal3 ;
  RECT 3094.480 0.000 3095.600 1.120 ;
  LAYER metal2 ;
  RECT 3094.480 0.000 3095.600 1.120 ;
  LAYER metal1 ;
  RECT 3094.480 0.000 3095.600 1.120 ;
 END
END DIA111
PIN DOA111
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3080.840 0.000 3081.960 1.120 ;
  LAYER metal4 ;
  RECT 3080.840 0.000 3081.960 1.120 ;
  LAYER metal3 ;
  RECT 3080.840 0.000 3081.960 1.120 ;
  LAYER metal2 ;
  RECT 3080.840 0.000 3081.960 1.120 ;
  LAYER metal1 ;
  RECT 3080.840 0.000 3081.960 1.120 ;
 END
END DOA111
PIN DIA110
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3067.820 0.000 3068.940 1.120 ;
  LAYER metal4 ;
  RECT 3067.820 0.000 3068.940 1.120 ;
  LAYER metal3 ;
  RECT 3067.820 0.000 3068.940 1.120 ;
  LAYER metal2 ;
  RECT 3067.820 0.000 3068.940 1.120 ;
  LAYER metal1 ;
  RECT 3067.820 0.000 3068.940 1.120 ;
 END
END DIA110
PIN DOA110
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3054.180 0.000 3055.300 1.120 ;
  LAYER metal4 ;
  RECT 3054.180 0.000 3055.300 1.120 ;
  LAYER metal3 ;
  RECT 3054.180 0.000 3055.300 1.120 ;
  LAYER metal2 ;
  RECT 3054.180 0.000 3055.300 1.120 ;
  LAYER metal1 ;
  RECT 3054.180 0.000 3055.300 1.120 ;
 END
END DOA110
PIN DIA109
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3040.540 0.000 3041.660 1.120 ;
  LAYER metal4 ;
  RECT 3040.540 0.000 3041.660 1.120 ;
  LAYER metal3 ;
  RECT 3040.540 0.000 3041.660 1.120 ;
  LAYER metal2 ;
  RECT 3040.540 0.000 3041.660 1.120 ;
  LAYER metal1 ;
  RECT 3040.540 0.000 3041.660 1.120 ;
 END
END DIA109
PIN DOA109
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3027.520 0.000 3028.640 1.120 ;
  LAYER metal4 ;
  RECT 3027.520 0.000 3028.640 1.120 ;
  LAYER metal3 ;
  RECT 3027.520 0.000 3028.640 1.120 ;
  LAYER metal2 ;
  RECT 3027.520 0.000 3028.640 1.120 ;
  LAYER metal1 ;
  RECT 3027.520 0.000 3028.640 1.120 ;
 END
END DOA109
PIN DIA108
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3013.880 0.000 3015.000 1.120 ;
  LAYER metal4 ;
  RECT 3013.880 0.000 3015.000 1.120 ;
  LAYER metal3 ;
  RECT 3013.880 0.000 3015.000 1.120 ;
  LAYER metal2 ;
  RECT 3013.880 0.000 3015.000 1.120 ;
  LAYER metal1 ;
  RECT 3013.880 0.000 3015.000 1.120 ;
 END
END DIA108
PIN DOA108
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3000.240 0.000 3001.360 1.120 ;
  LAYER metal4 ;
  RECT 3000.240 0.000 3001.360 1.120 ;
  LAYER metal3 ;
  RECT 3000.240 0.000 3001.360 1.120 ;
  LAYER metal2 ;
  RECT 3000.240 0.000 3001.360 1.120 ;
  LAYER metal1 ;
  RECT 3000.240 0.000 3001.360 1.120 ;
 END
END DOA108
PIN DIA107
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2987.220 0.000 2988.340 1.120 ;
  LAYER metal4 ;
  RECT 2987.220 0.000 2988.340 1.120 ;
  LAYER metal3 ;
  RECT 2987.220 0.000 2988.340 1.120 ;
  LAYER metal2 ;
  RECT 2987.220 0.000 2988.340 1.120 ;
  LAYER metal1 ;
  RECT 2987.220 0.000 2988.340 1.120 ;
 END
END DIA107
PIN DOA107
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2973.580 0.000 2974.700 1.120 ;
  LAYER metal4 ;
  RECT 2973.580 0.000 2974.700 1.120 ;
  LAYER metal3 ;
  RECT 2973.580 0.000 2974.700 1.120 ;
  LAYER metal2 ;
  RECT 2973.580 0.000 2974.700 1.120 ;
  LAYER metal1 ;
  RECT 2973.580 0.000 2974.700 1.120 ;
 END
END DOA107
PIN DIA106
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2959.940 0.000 2961.060 1.120 ;
  LAYER metal4 ;
  RECT 2959.940 0.000 2961.060 1.120 ;
  LAYER metal3 ;
  RECT 2959.940 0.000 2961.060 1.120 ;
  LAYER metal2 ;
  RECT 2959.940 0.000 2961.060 1.120 ;
  LAYER metal1 ;
  RECT 2959.940 0.000 2961.060 1.120 ;
 END
END DIA106
PIN DOA106
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2946.920 0.000 2948.040 1.120 ;
  LAYER metal4 ;
  RECT 2946.920 0.000 2948.040 1.120 ;
  LAYER metal3 ;
  RECT 2946.920 0.000 2948.040 1.120 ;
  LAYER metal2 ;
  RECT 2946.920 0.000 2948.040 1.120 ;
  LAYER metal1 ;
  RECT 2946.920 0.000 2948.040 1.120 ;
 END
END DOA106
PIN DIA105
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2933.280 0.000 2934.400 1.120 ;
  LAYER metal4 ;
  RECT 2933.280 0.000 2934.400 1.120 ;
  LAYER metal3 ;
  RECT 2933.280 0.000 2934.400 1.120 ;
  LAYER metal2 ;
  RECT 2933.280 0.000 2934.400 1.120 ;
  LAYER metal1 ;
  RECT 2933.280 0.000 2934.400 1.120 ;
 END
END DIA105
PIN DOA105
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2919.640 0.000 2920.760 1.120 ;
  LAYER metal4 ;
  RECT 2919.640 0.000 2920.760 1.120 ;
  LAYER metal3 ;
  RECT 2919.640 0.000 2920.760 1.120 ;
  LAYER metal2 ;
  RECT 2919.640 0.000 2920.760 1.120 ;
  LAYER metal1 ;
  RECT 2919.640 0.000 2920.760 1.120 ;
 END
END DOA105
PIN DIA104
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2906.000 0.000 2907.120 1.120 ;
  LAYER metal4 ;
  RECT 2906.000 0.000 2907.120 1.120 ;
  LAYER metal3 ;
  RECT 2906.000 0.000 2907.120 1.120 ;
  LAYER metal2 ;
  RECT 2906.000 0.000 2907.120 1.120 ;
  LAYER metal1 ;
  RECT 2906.000 0.000 2907.120 1.120 ;
 END
END DIA104
PIN DOA104
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2892.980 0.000 2894.100 1.120 ;
  LAYER metal4 ;
  RECT 2892.980 0.000 2894.100 1.120 ;
  LAYER metal3 ;
  RECT 2892.980 0.000 2894.100 1.120 ;
  LAYER metal2 ;
  RECT 2892.980 0.000 2894.100 1.120 ;
  LAYER metal1 ;
  RECT 2892.980 0.000 2894.100 1.120 ;
 END
END DOA104
PIN DIA103
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2879.340 0.000 2880.460 1.120 ;
  LAYER metal4 ;
  RECT 2879.340 0.000 2880.460 1.120 ;
  LAYER metal3 ;
  RECT 2879.340 0.000 2880.460 1.120 ;
  LAYER metal2 ;
  RECT 2879.340 0.000 2880.460 1.120 ;
  LAYER metal1 ;
  RECT 2879.340 0.000 2880.460 1.120 ;
 END
END DIA103
PIN DOA103
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2865.700 0.000 2866.820 1.120 ;
  LAYER metal4 ;
  RECT 2865.700 0.000 2866.820 1.120 ;
  LAYER metal3 ;
  RECT 2865.700 0.000 2866.820 1.120 ;
  LAYER metal2 ;
  RECT 2865.700 0.000 2866.820 1.120 ;
  LAYER metal1 ;
  RECT 2865.700 0.000 2866.820 1.120 ;
 END
END DOA103
PIN DIA102
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2852.680 0.000 2853.800 1.120 ;
  LAYER metal4 ;
  RECT 2852.680 0.000 2853.800 1.120 ;
  LAYER metal3 ;
  RECT 2852.680 0.000 2853.800 1.120 ;
  LAYER metal2 ;
  RECT 2852.680 0.000 2853.800 1.120 ;
  LAYER metal1 ;
  RECT 2852.680 0.000 2853.800 1.120 ;
 END
END DIA102
PIN DOA102
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2839.040 0.000 2840.160 1.120 ;
  LAYER metal4 ;
  RECT 2839.040 0.000 2840.160 1.120 ;
  LAYER metal3 ;
  RECT 2839.040 0.000 2840.160 1.120 ;
  LAYER metal2 ;
  RECT 2839.040 0.000 2840.160 1.120 ;
  LAYER metal1 ;
  RECT 2839.040 0.000 2840.160 1.120 ;
 END
END DOA102
PIN DIA101
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2825.400 0.000 2826.520 1.120 ;
  LAYER metal4 ;
  RECT 2825.400 0.000 2826.520 1.120 ;
  LAYER metal3 ;
  RECT 2825.400 0.000 2826.520 1.120 ;
  LAYER metal2 ;
  RECT 2825.400 0.000 2826.520 1.120 ;
  LAYER metal1 ;
  RECT 2825.400 0.000 2826.520 1.120 ;
 END
END DIA101
PIN DOA101
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2812.380 0.000 2813.500 1.120 ;
  LAYER metal4 ;
  RECT 2812.380 0.000 2813.500 1.120 ;
  LAYER metal3 ;
  RECT 2812.380 0.000 2813.500 1.120 ;
  LAYER metal2 ;
  RECT 2812.380 0.000 2813.500 1.120 ;
  LAYER metal1 ;
  RECT 2812.380 0.000 2813.500 1.120 ;
 END
END DOA101
PIN DIA100
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2798.740 0.000 2799.860 1.120 ;
  LAYER metal4 ;
  RECT 2798.740 0.000 2799.860 1.120 ;
  LAYER metal3 ;
  RECT 2798.740 0.000 2799.860 1.120 ;
  LAYER metal2 ;
  RECT 2798.740 0.000 2799.860 1.120 ;
  LAYER metal1 ;
  RECT 2798.740 0.000 2799.860 1.120 ;
 END
END DIA100
PIN DOA100
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2785.100 0.000 2786.220 1.120 ;
  LAYER metal4 ;
  RECT 2785.100 0.000 2786.220 1.120 ;
  LAYER metal3 ;
  RECT 2785.100 0.000 2786.220 1.120 ;
  LAYER metal2 ;
  RECT 2785.100 0.000 2786.220 1.120 ;
  LAYER metal1 ;
  RECT 2785.100 0.000 2786.220 1.120 ;
 END
END DOA100
PIN DIA99
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2772.080 0.000 2773.200 1.120 ;
  LAYER metal4 ;
  RECT 2772.080 0.000 2773.200 1.120 ;
  LAYER metal3 ;
  RECT 2772.080 0.000 2773.200 1.120 ;
  LAYER metal2 ;
  RECT 2772.080 0.000 2773.200 1.120 ;
  LAYER metal1 ;
  RECT 2772.080 0.000 2773.200 1.120 ;
 END
END DIA99
PIN DOA99
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2758.440 0.000 2759.560 1.120 ;
  LAYER metal4 ;
  RECT 2758.440 0.000 2759.560 1.120 ;
  LAYER metal3 ;
  RECT 2758.440 0.000 2759.560 1.120 ;
  LAYER metal2 ;
  RECT 2758.440 0.000 2759.560 1.120 ;
  LAYER metal1 ;
  RECT 2758.440 0.000 2759.560 1.120 ;
 END
END DOA99
PIN DIA98
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2744.800 0.000 2745.920 1.120 ;
  LAYER metal4 ;
  RECT 2744.800 0.000 2745.920 1.120 ;
  LAYER metal3 ;
  RECT 2744.800 0.000 2745.920 1.120 ;
  LAYER metal2 ;
  RECT 2744.800 0.000 2745.920 1.120 ;
  LAYER metal1 ;
  RECT 2744.800 0.000 2745.920 1.120 ;
 END
END DIA98
PIN DOA98
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2731.780 0.000 2732.900 1.120 ;
  LAYER metal4 ;
  RECT 2731.780 0.000 2732.900 1.120 ;
  LAYER metal3 ;
  RECT 2731.780 0.000 2732.900 1.120 ;
  LAYER metal2 ;
  RECT 2731.780 0.000 2732.900 1.120 ;
  LAYER metal1 ;
  RECT 2731.780 0.000 2732.900 1.120 ;
 END
END DOA98
PIN DIA97
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2718.140 0.000 2719.260 1.120 ;
  LAYER metal4 ;
  RECT 2718.140 0.000 2719.260 1.120 ;
  LAYER metal3 ;
  RECT 2718.140 0.000 2719.260 1.120 ;
  LAYER metal2 ;
  RECT 2718.140 0.000 2719.260 1.120 ;
  LAYER metal1 ;
  RECT 2718.140 0.000 2719.260 1.120 ;
 END
END DIA97
PIN DOA97
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2704.500 0.000 2705.620 1.120 ;
  LAYER metal4 ;
  RECT 2704.500 0.000 2705.620 1.120 ;
  LAYER metal3 ;
  RECT 2704.500 0.000 2705.620 1.120 ;
  LAYER metal2 ;
  RECT 2704.500 0.000 2705.620 1.120 ;
  LAYER metal1 ;
  RECT 2704.500 0.000 2705.620 1.120 ;
 END
END DOA97
PIN DIA96
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2691.480 0.000 2692.600 1.120 ;
  LAYER metal4 ;
  RECT 2691.480 0.000 2692.600 1.120 ;
  LAYER metal3 ;
  RECT 2691.480 0.000 2692.600 1.120 ;
  LAYER metal2 ;
  RECT 2691.480 0.000 2692.600 1.120 ;
  LAYER metal1 ;
  RECT 2691.480 0.000 2692.600 1.120 ;
 END
END DIA96
PIN WEAN6
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 2680.320 0.000 2681.440 1.120 ;
  LAYER metal4 ;
  RECT 2680.320 0.000 2681.440 1.120 ;
  LAYER metal3 ;
  RECT 2680.320 0.000 2681.440 1.120 ;
  LAYER metal2 ;
  RECT 2680.320 0.000 2681.440 1.120 ;
  LAYER metal1 ;
  RECT 2680.320 0.000 2681.440 1.120 ;
 END
END WEAN6
PIN DOA96
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2677.840 0.000 2678.960 1.120 ;
  LAYER metal4 ;
  RECT 2677.840 0.000 2678.960 1.120 ;
  LAYER metal3 ;
  RECT 2677.840 0.000 2678.960 1.120 ;
  LAYER metal2 ;
  RECT 2677.840 0.000 2678.960 1.120 ;
  LAYER metal1 ;
  RECT 2677.840 0.000 2678.960 1.120 ;
 END
END DOA96
PIN DIA95
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2664.200 0.000 2665.320 1.120 ;
  LAYER metal4 ;
  RECT 2664.200 0.000 2665.320 1.120 ;
  LAYER metal3 ;
  RECT 2664.200 0.000 2665.320 1.120 ;
  LAYER metal2 ;
  RECT 2664.200 0.000 2665.320 1.120 ;
  LAYER metal1 ;
  RECT 2664.200 0.000 2665.320 1.120 ;
 END
END DIA95
PIN DOA95
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2651.180 0.000 2652.300 1.120 ;
  LAYER metal4 ;
  RECT 2651.180 0.000 2652.300 1.120 ;
  LAYER metal3 ;
  RECT 2651.180 0.000 2652.300 1.120 ;
  LAYER metal2 ;
  RECT 2651.180 0.000 2652.300 1.120 ;
  LAYER metal1 ;
  RECT 2651.180 0.000 2652.300 1.120 ;
 END
END DOA95
PIN DIA94
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2637.540 0.000 2638.660 1.120 ;
  LAYER metal4 ;
  RECT 2637.540 0.000 2638.660 1.120 ;
  LAYER metal3 ;
  RECT 2637.540 0.000 2638.660 1.120 ;
  LAYER metal2 ;
  RECT 2637.540 0.000 2638.660 1.120 ;
  LAYER metal1 ;
  RECT 2637.540 0.000 2638.660 1.120 ;
 END
END DIA94
PIN DOA94
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2623.900 0.000 2625.020 1.120 ;
  LAYER metal4 ;
  RECT 2623.900 0.000 2625.020 1.120 ;
  LAYER metal3 ;
  RECT 2623.900 0.000 2625.020 1.120 ;
  LAYER metal2 ;
  RECT 2623.900 0.000 2625.020 1.120 ;
  LAYER metal1 ;
  RECT 2623.900 0.000 2625.020 1.120 ;
 END
END DOA94
PIN DIA93
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2610.880 0.000 2612.000 1.120 ;
  LAYER metal4 ;
  RECT 2610.880 0.000 2612.000 1.120 ;
  LAYER metal3 ;
  RECT 2610.880 0.000 2612.000 1.120 ;
  LAYER metal2 ;
  RECT 2610.880 0.000 2612.000 1.120 ;
  LAYER metal1 ;
  RECT 2610.880 0.000 2612.000 1.120 ;
 END
END DIA93
PIN DOA93
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2597.240 0.000 2598.360 1.120 ;
  LAYER metal4 ;
  RECT 2597.240 0.000 2598.360 1.120 ;
  LAYER metal3 ;
  RECT 2597.240 0.000 2598.360 1.120 ;
  LAYER metal2 ;
  RECT 2597.240 0.000 2598.360 1.120 ;
  LAYER metal1 ;
  RECT 2597.240 0.000 2598.360 1.120 ;
 END
END DOA93
PIN DIA92
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2583.600 0.000 2584.720 1.120 ;
  LAYER metal4 ;
  RECT 2583.600 0.000 2584.720 1.120 ;
  LAYER metal3 ;
  RECT 2583.600 0.000 2584.720 1.120 ;
  LAYER metal2 ;
  RECT 2583.600 0.000 2584.720 1.120 ;
  LAYER metal1 ;
  RECT 2583.600 0.000 2584.720 1.120 ;
 END
END DIA92
PIN DOA92
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2570.580 0.000 2571.700 1.120 ;
  LAYER metal4 ;
  RECT 2570.580 0.000 2571.700 1.120 ;
  LAYER metal3 ;
  RECT 2570.580 0.000 2571.700 1.120 ;
  LAYER metal2 ;
  RECT 2570.580 0.000 2571.700 1.120 ;
  LAYER metal1 ;
  RECT 2570.580 0.000 2571.700 1.120 ;
 END
END DOA92
PIN DIA91
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2556.940 0.000 2558.060 1.120 ;
  LAYER metal4 ;
  RECT 2556.940 0.000 2558.060 1.120 ;
  LAYER metal3 ;
  RECT 2556.940 0.000 2558.060 1.120 ;
  LAYER metal2 ;
  RECT 2556.940 0.000 2558.060 1.120 ;
  LAYER metal1 ;
  RECT 2556.940 0.000 2558.060 1.120 ;
 END
END DIA91
PIN DOA91
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2543.300 0.000 2544.420 1.120 ;
  LAYER metal4 ;
  RECT 2543.300 0.000 2544.420 1.120 ;
  LAYER metal3 ;
  RECT 2543.300 0.000 2544.420 1.120 ;
  LAYER metal2 ;
  RECT 2543.300 0.000 2544.420 1.120 ;
  LAYER metal1 ;
  RECT 2543.300 0.000 2544.420 1.120 ;
 END
END DOA91
PIN DIA90
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2530.280 0.000 2531.400 1.120 ;
  LAYER metal4 ;
  RECT 2530.280 0.000 2531.400 1.120 ;
  LAYER metal3 ;
  RECT 2530.280 0.000 2531.400 1.120 ;
  LAYER metal2 ;
  RECT 2530.280 0.000 2531.400 1.120 ;
  LAYER metal1 ;
  RECT 2530.280 0.000 2531.400 1.120 ;
 END
END DIA90
PIN DOA90
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2516.640 0.000 2517.760 1.120 ;
  LAYER metal4 ;
  RECT 2516.640 0.000 2517.760 1.120 ;
  LAYER metal3 ;
  RECT 2516.640 0.000 2517.760 1.120 ;
  LAYER metal2 ;
  RECT 2516.640 0.000 2517.760 1.120 ;
  LAYER metal1 ;
  RECT 2516.640 0.000 2517.760 1.120 ;
 END
END DOA90
PIN DIA89
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2503.000 0.000 2504.120 1.120 ;
  LAYER metal4 ;
  RECT 2503.000 0.000 2504.120 1.120 ;
  LAYER metal3 ;
  RECT 2503.000 0.000 2504.120 1.120 ;
  LAYER metal2 ;
  RECT 2503.000 0.000 2504.120 1.120 ;
  LAYER metal1 ;
  RECT 2503.000 0.000 2504.120 1.120 ;
 END
END DIA89
PIN DOA89
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2489.360 0.000 2490.480 1.120 ;
  LAYER metal4 ;
  RECT 2489.360 0.000 2490.480 1.120 ;
  LAYER metal3 ;
  RECT 2489.360 0.000 2490.480 1.120 ;
  LAYER metal2 ;
  RECT 2489.360 0.000 2490.480 1.120 ;
  LAYER metal1 ;
  RECT 2489.360 0.000 2490.480 1.120 ;
 END
END DOA89
PIN DIA88
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2476.340 0.000 2477.460 1.120 ;
  LAYER metal4 ;
  RECT 2476.340 0.000 2477.460 1.120 ;
  LAYER metal3 ;
  RECT 2476.340 0.000 2477.460 1.120 ;
  LAYER metal2 ;
  RECT 2476.340 0.000 2477.460 1.120 ;
  LAYER metal1 ;
  RECT 2476.340 0.000 2477.460 1.120 ;
 END
END DIA88
PIN DOA88
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2462.700 0.000 2463.820 1.120 ;
  LAYER metal4 ;
  RECT 2462.700 0.000 2463.820 1.120 ;
  LAYER metal3 ;
  RECT 2462.700 0.000 2463.820 1.120 ;
  LAYER metal2 ;
  RECT 2462.700 0.000 2463.820 1.120 ;
  LAYER metal1 ;
  RECT 2462.700 0.000 2463.820 1.120 ;
 END
END DOA88
PIN DIA87
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2449.060 0.000 2450.180 1.120 ;
  LAYER metal4 ;
  RECT 2449.060 0.000 2450.180 1.120 ;
  LAYER metal3 ;
  RECT 2449.060 0.000 2450.180 1.120 ;
  LAYER metal2 ;
  RECT 2449.060 0.000 2450.180 1.120 ;
  LAYER metal1 ;
  RECT 2449.060 0.000 2450.180 1.120 ;
 END
END DIA87
PIN DOA87
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2436.040 0.000 2437.160 1.120 ;
  LAYER metal4 ;
  RECT 2436.040 0.000 2437.160 1.120 ;
  LAYER metal3 ;
  RECT 2436.040 0.000 2437.160 1.120 ;
  LAYER metal2 ;
  RECT 2436.040 0.000 2437.160 1.120 ;
  LAYER metal1 ;
  RECT 2436.040 0.000 2437.160 1.120 ;
 END
END DOA87
PIN DIA86
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2422.400 0.000 2423.520 1.120 ;
  LAYER metal4 ;
  RECT 2422.400 0.000 2423.520 1.120 ;
  LAYER metal3 ;
  RECT 2422.400 0.000 2423.520 1.120 ;
  LAYER metal2 ;
  RECT 2422.400 0.000 2423.520 1.120 ;
  LAYER metal1 ;
  RECT 2422.400 0.000 2423.520 1.120 ;
 END
END DIA86
PIN DOA86
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2408.760 0.000 2409.880 1.120 ;
  LAYER metal4 ;
  RECT 2408.760 0.000 2409.880 1.120 ;
  LAYER metal3 ;
  RECT 2408.760 0.000 2409.880 1.120 ;
  LAYER metal2 ;
  RECT 2408.760 0.000 2409.880 1.120 ;
  LAYER metal1 ;
  RECT 2408.760 0.000 2409.880 1.120 ;
 END
END DOA86
PIN DIA85
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2395.740 0.000 2396.860 1.120 ;
  LAYER metal4 ;
  RECT 2395.740 0.000 2396.860 1.120 ;
  LAYER metal3 ;
  RECT 2395.740 0.000 2396.860 1.120 ;
  LAYER metal2 ;
  RECT 2395.740 0.000 2396.860 1.120 ;
  LAYER metal1 ;
  RECT 2395.740 0.000 2396.860 1.120 ;
 END
END DIA85
PIN DOA85
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2382.100 0.000 2383.220 1.120 ;
  LAYER metal4 ;
  RECT 2382.100 0.000 2383.220 1.120 ;
  LAYER metal3 ;
  RECT 2382.100 0.000 2383.220 1.120 ;
  LAYER metal2 ;
  RECT 2382.100 0.000 2383.220 1.120 ;
  LAYER metal1 ;
  RECT 2382.100 0.000 2383.220 1.120 ;
 END
END DOA85
PIN DIA84
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2368.460 0.000 2369.580 1.120 ;
  LAYER metal4 ;
  RECT 2368.460 0.000 2369.580 1.120 ;
  LAYER metal3 ;
  RECT 2368.460 0.000 2369.580 1.120 ;
  LAYER metal2 ;
  RECT 2368.460 0.000 2369.580 1.120 ;
  LAYER metal1 ;
  RECT 2368.460 0.000 2369.580 1.120 ;
 END
END DIA84
PIN DOA84
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2355.440 0.000 2356.560 1.120 ;
  LAYER metal4 ;
  RECT 2355.440 0.000 2356.560 1.120 ;
  LAYER metal3 ;
  RECT 2355.440 0.000 2356.560 1.120 ;
  LAYER metal2 ;
  RECT 2355.440 0.000 2356.560 1.120 ;
  LAYER metal1 ;
  RECT 2355.440 0.000 2356.560 1.120 ;
 END
END DOA84
PIN DIA83
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2341.800 0.000 2342.920 1.120 ;
  LAYER metal4 ;
  RECT 2341.800 0.000 2342.920 1.120 ;
  LAYER metal3 ;
  RECT 2341.800 0.000 2342.920 1.120 ;
  LAYER metal2 ;
  RECT 2341.800 0.000 2342.920 1.120 ;
  LAYER metal1 ;
  RECT 2341.800 0.000 2342.920 1.120 ;
 END
END DIA83
PIN DOA83
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2328.160 0.000 2329.280 1.120 ;
  LAYER metal4 ;
  RECT 2328.160 0.000 2329.280 1.120 ;
  LAYER metal3 ;
  RECT 2328.160 0.000 2329.280 1.120 ;
  LAYER metal2 ;
  RECT 2328.160 0.000 2329.280 1.120 ;
  LAYER metal1 ;
  RECT 2328.160 0.000 2329.280 1.120 ;
 END
END DOA83
PIN DIA82
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2315.140 0.000 2316.260 1.120 ;
  LAYER metal4 ;
  RECT 2315.140 0.000 2316.260 1.120 ;
  LAYER metal3 ;
  RECT 2315.140 0.000 2316.260 1.120 ;
  LAYER metal2 ;
  RECT 2315.140 0.000 2316.260 1.120 ;
  LAYER metal1 ;
  RECT 2315.140 0.000 2316.260 1.120 ;
 END
END DIA82
PIN DOA82
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2301.500 0.000 2302.620 1.120 ;
  LAYER metal4 ;
  RECT 2301.500 0.000 2302.620 1.120 ;
  LAYER metal3 ;
  RECT 2301.500 0.000 2302.620 1.120 ;
  LAYER metal2 ;
  RECT 2301.500 0.000 2302.620 1.120 ;
  LAYER metal1 ;
  RECT 2301.500 0.000 2302.620 1.120 ;
 END
END DOA82
PIN DIA81
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2287.860 0.000 2288.980 1.120 ;
  LAYER metal4 ;
  RECT 2287.860 0.000 2288.980 1.120 ;
  LAYER metal3 ;
  RECT 2287.860 0.000 2288.980 1.120 ;
  LAYER metal2 ;
  RECT 2287.860 0.000 2288.980 1.120 ;
  LAYER metal1 ;
  RECT 2287.860 0.000 2288.980 1.120 ;
 END
END DIA81
PIN DOA81
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2274.840 0.000 2275.960 1.120 ;
  LAYER metal4 ;
  RECT 2274.840 0.000 2275.960 1.120 ;
  LAYER metal3 ;
  RECT 2274.840 0.000 2275.960 1.120 ;
  LAYER metal2 ;
  RECT 2274.840 0.000 2275.960 1.120 ;
  LAYER metal1 ;
  RECT 2274.840 0.000 2275.960 1.120 ;
 END
END DOA81
PIN DIA80
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2261.200 0.000 2262.320 1.120 ;
  LAYER metal4 ;
  RECT 2261.200 0.000 2262.320 1.120 ;
  LAYER metal3 ;
  RECT 2261.200 0.000 2262.320 1.120 ;
  LAYER metal2 ;
  RECT 2261.200 0.000 2262.320 1.120 ;
  LAYER metal1 ;
  RECT 2261.200 0.000 2262.320 1.120 ;
 END
END DIA80
PIN WEAN5
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 2250.040 0.000 2251.160 1.120 ;
  LAYER metal4 ;
  RECT 2250.040 0.000 2251.160 1.120 ;
  LAYER metal3 ;
  RECT 2250.040 0.000 2251.160 1.120 ;
  LAYER metal2 ;
  RECT 2250.040 0.000 2251.160 1.120 ;
  LAYER metal1 ;
  RECT 2250.040 0.000 2251.160 1.120 ;
 END
END WEAN5
PIN DOA80
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2247.560 0.000 2248.680 1.120 ;
  LAYER metal4 ;
  RECT 2247.560 0.000 2248.680 1.120 ;
  LAYER metal3 ;
  RECT 2247.560 0.000 2248.680 1.120 ;
  LAYER metal2 ;
  RECT 2247.560 0.000 2248.680 1.120 ;
  LAYER metal1 ;
  RECT 2247.560 0.000 2248.680 1.120 ;
 END
END DOA80
PIN DIA79
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2234.540 0.000 2235.660 1.120 ;
  LAYER metal4 ;
  RECT 2234.540 0.000 2235.660 1.120 ;
  LAYER metal3 ;
  RECT 2234.540 0.000 2235.660 1.120 ;
  LAYER metal2 ;
  RECT 2234.540 0.000 2235.660 1.120 ;
  LAYER metal1 ;
  RECT 2234.540 0.000 2235.660 1.120 ;
 END
END DIA79
PIN DOA79
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2220.900 0.000 2222.020 1.120 ;
  LAYER metal4 ;
  RECT 2220.900 0.000 2222.020 1.120 ;
  LAYER metal3 ;
  RECT 2220.900 0.000 2222.020 1.120 ;
  LAYER metal2 ;
  RECT 2220.900 0.000 2222.020 1.120 ;
  LAYER metal1 ;
  RECT 2220.900 0.000 2222.020 1.120 ;
 END
END DOA79
PIN DIA78
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2207.260 0.000 2208.380 1.120 ;
  LAYER metal4 ;
  RECT 2207.260 0.000 2208.380 1.120 ;
  LAYER metal3 ;
  RECT 2207.260 0.000 2208.380 1.120 ;
  LAYER metal2 ;
  RECT 2207.260 0.000 2208.380 1.120 ;
  LAYER metal1 ;
  RECT 2207.260 0.000 2208.380 1.120 ;
 END
END DIA78
PIN DOA78
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2194.240 0.000 2195.360 1.120 ;
  LAYER metal4 ;
  RECT 2194.240 0.000 2195.360 1.120 ;
  LAYER metal3 ;
  RECT 2194.240 0.000 2195.360 1.120 ;
  LAYER metal2 ;
  RECT 2194.240 0.000 2195.360 1.120 ;
  LAYER metal1 ;
  RECT 2194.240 0.000 2195.360 1.120 ;
 END
END DOA78
PIN DIA77
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2180.600 0.000 2181.720 1.120 ;
  LAYER metal4 ;
  RECT 2180.600 0.000 2181.720 1.120 ;
  LAYER metal3 ;
  RECT 2180.600 0.000 2181.720 1.120 ;
  LAYER metal2 ;
  RECT 2180.600 0.000 2181.720 1.120 ;
  LAYER metal1 ;
  RECT 2180.600 0.000 2181.720 1.120 ;
 END
END DIA77
PIN DOA77
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2166.960 0.000 2168.080 1.120 ;
  LAYER metal4 ;
  RECT 2166.960 0.000 2168.080 1.120 ;
  LAYER metal3 ;
  RECT 2166.960 0.000 2168.080 1.120 ;
  LAYER metal2 ;
  RECT 2166.960 0.000 2168.080 1.120 ;
  LAYER metal1 ;
  RECT 2166.960 0.000 2168.080 1.120 ;
 END
END DOA77
PIN DIA76
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2153.940 0.000 2155.060 1.120 ;
  LAYER metal4 ;
  RECT 2153.940 0.000 2155.060 1.120 ;
  LAYER metal3 ;
  RECT 2153.940 0.000 2155.060 1.120 ;
  LAYER metal2 ;
  RECT 2153.940 0.000 2155.060 1.120 ;
  LAYER metal1 ;
  RECT 2153.940 0.000 2155.060 1.120 ;
 END
END DIA76
PIN DOA76
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2140.300 0.000 2141.420 1.120 ;
  LAYER metal4 ;
  RECT 2140.300 0.000 2141.420 1.120 ;
  LAYER metal3 ;
  RECT 2140.300 0.000 2141.420 1.120 ;
  LAYER metal2 ;
  RECT 2140.300 0.000 2141.420 1.120 ;
  LAYER metal1 ;
  RECT 2140.300 0.000 2141.420 1.120 ;
 END
END DOA76
PIN DIA75
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2126.660 0.000 2127.780 1.120 ;
  LAYER metal4 ;
  RECT 2126.660 0.000 2127.780 1.120 ;
  LAYER metal3 ;
  RECT 2126.660 0.000 2127.780 1.120 ;
  LAYER metal2 ;
  RECT 2126.660 0.000 2127.780 1.120 ;
  LAYER metal1 ;
  RECT 2126.660 0.000 2127.780 1.120 ;
 END
END DIA75
PIN DOA75
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2113.640 0.000 2114.760 1.120 ;
  LAYER metal4 ;
  RECT 2113.640 0.000 2114.760 1.120 ;
  LAYER metal3 ;
  RECT 2113.640 0.000 2114.760 1.120 ;
  LAYER metal2 ;
  RECT 2113.640 0.000 2114.760 1.120 ;
  LAYER metal1 ;
  RECT 2113.640 0.000 2114.760 1.120 ;
 END
END DOA75
PIN DIA74
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2100.000 0.000 2101.120 1.120 ;
  LAYER metal4 ;
  RECT 2100.000 0.000 2101.120 1.120 ;
  LAYER metal3 ;
  RECT 2100.000 0.000 2101.120 1.120 ;
  LAYER metal2 ;
  RECT 2100.000 0.000 2101.120 1.120 ;
  LAYER metal1 ;
  RECT 2100.000 0.000 2101.120 1.120 ;
 END
END DIA74
PIN DOA74
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2086.360 0.000 2087.480 1.120 ;
  LAYER metal4 ;
  RECT 2086.360 0.000 2087.480 1.120 ;
  LAYER metal3 ;
  RECT 2086.360 0.000 2087.480 1.120 ;
  LAYER metal2 ;
  RECT 2086.360 0.000 2087.480 1.120 ;
  LAYER metal1 ;
  RECT 2086.360 0.000 2087.480 1.120 ;
 END
END DOA74
PIN DIA73
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2072.720 0.000 2073.840 1.120 ;
  LAYER metal4 ;
  RECT 2072.720 0.000 2073.840 1.120 ;
  LAYER metal3 ;
  RECT 2072.720 0.000 2073.840 1.120 ;
  LAYER metal2 ;
  RECT 2072.720 0.000 2073.840 1.120 ;
  LAYER metal1 ;
  RECT 2072.720 0.000 2073.840 1.120 ;
 END
END DIA73
PIN DOA73
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2059.700 0.000 2060.820 1.120 ;
  LAYER metal4 ;
  RECT 2059.700 0.000 2060.820 1.120 ;
  LAYER metal3 ;
  RECT 2059.700 0.000 2060.820 1.120 ;
  LAYER metal2 ;
  RECT 2059.700 0.000 2060.820 1.120 ;
  LAYER metal1 ;
  RECT 2059.700 0.000 2060.820 1.120 ;
 END
END DOA73
PIN DIA72
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2046.060 0.000 2047.180 1.120 ;
  LAYER metal4 ;
  RECT 2046.060 0.000 2047.180 1.120 ;
  LAYER metal3 ;
  RECT 2046.060 0.000 2047.180 1.120 ;
  LAYER metal2 ;
  RECT 2046.060 0.000 2047.180 1.120 ;
  LAYER metal1 ;
  RECT 2046.060 0.000 2047.180 1.120 ;
 END
END DIA72
PIN DOA72
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2032.420 0.000 2033.540 1.120 ;
  LAYER metal4 ;
  RECT 2032.420 0.000 2033.540 1.120 ;
  LAYER metal3 ;
  RECT 2032.420 0.000 2033.540 1.120 ;
  LAYER metal2 ;
  RECT 2032.420 0.000 2033.540 1.120 ;
  LAYER metal1 ;
  RECT 2032.420 0.000 2033.540 1.120 ;
 END
END DOA72
PIN DIA71
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2019.400 0.000 2020.520 1.120 ;
  LAYER metal4 ;
  RECT 2019.400 0.000 2020.520 1.120 ;
  LAYER metal3 ;
  RECT 2019.400 0.000 2020.520 1.120 ;
  LAYER metal2 ;
  RECT 2019.400 0.000 2020.520 1.120 ;
  LAYER metal1 ;
  RECT 2019.400 0.000 2020.520 1.120 ;
 END
END DIA71
PIN DOA71
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2005.760 0.000 2006.880 1.120 ;
  LAYER metal4 ;
  RECT 2005.760 0.000 2006.880 1.120 ;
  LAYER metal3 ;
  RECT 2005.760 0.000 2006.880 1.120 ;
  LAYER metal2 ;
  RECT 2005.760 0.000 2006.880 1.120 ;
  LAYER metal1 ;
  RECT 2005.760 0.000 2006.880 1.120 ;
 END
END DOA71
PIN DIA70
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1992.120 0.000 1993.240 1.120 ;
  LAYER metal4 ;
  RECT 1992.120 0.000 1993.240 1.120 ;
  LAYER metal3 ;
  RECT 1992.120 0.000 1993.240 1.120 ;
  LAYER metal2 ;
  RECT 1992.120 0.000 1993.240 1.120 ;
  LAYER metal1 ;
  RECT 1992.120 0.000 1993.240 1.120 ;
 END
END DIA70
PIN DOA70
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1979.100 0.000 1980.220 1.120 ;
  LAYER metal4 ;
  RECT 1979.100 0.000 1980.220 1.120 ;
  LAYER metal3 ;
  RECT 1979.100 0.000 1980.220 1.120 ;
  LAYER metal2 ;
  RECT 1979.100 0.000 1980.220 1.120 ;
  LAYER metal1 ;
  RECT 1979.100 0.000 1980.220 1.120 ;
 END
END DOA70
PIN DIA69
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1965.460 0.000 1966.580 1.120 ;
  LAYER metal4 ;
  RECT 1965.460 0.000 1966.580 1.120 ;
  LAYER metal3 ;
  RECT 1965.460 0.000 1966.580 1.120 ;
  LAYER metal2 ;
  RECT 1965.460 0.000 1966.580 1.120 ;
  LAYER metal1 ;
  RECT 1965.460 0.000 1966.580 1.120 ;
 END
END DIA69
PIN DOA69
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1951.820 0.000 1952.940 1.120 ;
  LAYER metal4 ;
  RECT 1951.820 0.000 1952.940 1.120 ;
  LAYER metal3 ;
  RECT 1951.820 0.000 1952.940 1.120 ;
  LAYER metal2 ;
  RECT 1951.820 0.000 1952.940 1.120 ;
  LAYER metal1 ;
  RECT 1951.820 0.000 1952.940 1.120 ;
 END
END DOA69
PIN DIA68
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1938.800 0.000 1939.920 1.120 ;
  LAYER metal4 ;
  RECT 1938.800 0.000 1939.920 1.120 ;
  LAYER metal3 ;
  RECT 1938.800 0.000 1939.920 1.120 ;
  LAYER metal2 ;
  RECT 1938.800 0.000 1939.920 1.120 ;
  LAYER metal1 ;
  RECT 1938.800 0.000 1939.920 1.120 ;
 END
END DIA68
PIN DOA68
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1925.160 0.000 1926.280 1.120 ;
  LAYER metal4 ;
  RECT 1925.160 0.000 1926.280 1.120 ;
  LAYER metal3 ;
  RECT 1925.160 0.000 1926.280 1.120 ;
  LAYER metal2 ;
  RECT 1925.160 0.000 1926.280 1.120 ;
  LAYER metal1 ;
  RECT 1925.160 0.000 1926.280 1.120 ;
 END
END DOA68
PIN DIA67
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1911.520 0.000 1912.640 1.120 ;
  LAYER metal4 ;
  RECT 1911.520 0.000 1912.640 1.120 ;
  LAYER metal3 ;
  RECT 1911.520 0.000 1912.640 1.120 ;
  LAYER metal2 ;
  RECT 1911.520 0.000 1912.640 1.120 ;
  LAYER metal1 ;
  RECT 1911.520 0.000 1912.640 1.120 ;
 END
END DIA67
PIN DOA67
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1898.500 0.000 1899.620 1.120 ;
  LAYER metal4 ;
  RECT 1898.500 0.000 1899.620 1.120 ;
  LAYER metal3 ;
  RECT 1898.500 0.000 1899.620 1.120 ;
  LAYER metal2 ;
  RECT 1898.500 0.000 1899.620 1.120 ;
  LAYER metal1 ;
  RECT 1898.500 0.000 1899.620 1.120 ;
 END
END DOA67
PIN DIA66
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1884.860 0.000 1885.980 1.120 ;
  LAYER metal4 ;
  RECT 1884.860 0.000 1885.980 1.120 ;
  LAYER metal3 ;
  RECT 1884.860 0.000 1885.980 1.120 ;
  LAYER metal2 ;
  RECT 1884.860 0.000 1885.980 1.120 ;
  LAYER metal1 ;
  RECT 1884.860 0.000 1885.980 1.120 ;
 END
END DIA66
PIN DOA66
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1871.220 0.000 1872.340 1.120 ;
  LAYER metal4 ;
  RECT 1871.220 0.000 1872.340 1.120 ;
  LAYER metal3 ;
  RECT 1871.220 0.000 1872.340 1.120 ;
  LAYER metal2 ;
  RECT 1871.220 0.000 1872.340 1.120 ;
  LAYER metal1 ;
  RECT 1871.220 0.000 1872.340 1.120 ;
 END
END DOA66
PIN DIA65
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1858.200 0.000 1859.320 1.120 ;
  LAYER metal4 ;
  RECT 1858.200 0.000 1859.320 1.120 ;
  LAYER metal3 ;
  RECT 1858.200 0.000 1859.320 1.120 ;
  LAYER metal2 ;
  RECT 1858.200 0.000 1859.320 1.120 ;
  LAYER metal1 ;
  RECT 1858.200 0.000 1859.320 1.120 ;
 END
END DIA65
PIN DOA65
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1844.560 0.000 1845.680 1.120 ;
  LAYER metal4 ;
  RECT 1844.560 0.000 1845.680 1.120 ;
  LAYER metal3 ;
  RECT 1844.560 0.000 1845.680 1.120 ;
  LAYER metal2 ;
  RECT 1844.560 0.000 1845.680 1.120 ;
  LAYER metal1 ;
  RECT 1844.560 0.000 1845.680 1.120 ;
 END
END DOA65
PIN DIA64
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1830.920 0.000 1832.040 1.120 ;
  LAYER metal4 ;
  RECT 1830.920 0.000 1832.040 1.120 ;
  LAYER metal3 ;
  RECT 1830.920 0.000 1832.040 1.120 ;
  LAYER metal2 ;
  RECT 1830.920 0.000 1832.040 1.120 ;
  LAYER metal1 ;
  RECT 1830.920 0.000 1832.040 1.120 ;
 END
END DIA64
PIN WEAN4
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1819.760 0.000 1820.880 1.120 ;
  LAYER metal4 ;
  RECT 1819.760 0.000 1820.880 1.120 ;
  LAYER metal3 ;
  RECT 1819.760 0.000 1820.880 1.120 ;
  LAYER metal2 ;
  RECT 1819.760 0.000 1820.880 1.120 ;
  LAYER metal1 ;
  RECT 1819.760 0.000 1820.880 1.120 ;
 END
END WEAN4
PIN DOA64
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1817.900 0.000 1819.020 1.120 ;
  LAYER metal4 ;
  RECT 1817.900 0.000 1819.020 1.120 ;
  LAYER metal3 ;
  RECT 1817.900 0.000 1819.020 1.120 ;
  LAYER metal2 ;
  RECT 1817.900 0.000 1819.020 1.120 ;
  LAYER metal1 ;
  RECT 1817.900 0.000 1819.020 1.120 ;
 END
END DOA64
PIN OEA
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1790.620 0.000 1791.740 1.120 ;
  LAYER metal4 ;
  RECT 1790.620 0.000 1791.740 1.120 ;
  LAYER metal3 ;
  RECT 1790.620 0.000 1791.740 1.120 ;
  LAYER metal2 ;
  RECT 1790.620 0.000 1791.740 1.120 ;
  LAYER metal1 ;
  RECT 1790.620 0.000 1791.740 1.120 ;
 END
END OEA
PIN CKA
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1777.600 0.000 1778.720 1.120 ;
  LAYER metal4 ;
  RECT 1777.600 0.000 1778.720 1.120 ;
  LAYER metal3 ;
  RECT 1777.600 0.000 1778.720 1.120 ;
  LAYER metal2 ;
  RECT 1777.600 0.000 1778.720 1.120 ;
  LAYER metal1 ;
  RECT 1777.600 0.000 1778.720 1.120 ;
 END
END CKA
PIN CSA
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1775.740 0.000 1776.860 1.120 ;
  LAYER metal4 ;
  RECT 1775.740 0.000 1776.860 1.120 ;
  LAYER metal3 ;
  RECT 1775.740 0.000 1776.860 1.120 ;
  LAYER metal2 ;
  RECT 1775.740 0.000 1776.860 1.120 ;
  LAYER metal1 ;
  RECT 1775.740 0.000 1776.860 1.120 ;
 END
END CSA
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1768.920 0.000 1770.040 1.120 ;
  LAYER metal4 ;
  RECT 1768.920 0.000 1770.040 1.120 ;
  LAYER metal3 ;
  RECT 1768.920 0.000 1770.040 1.120 ;
  LAYER metal2 ;
  RECT 1768.920 0.000 1770.040 1.120 ;
  LAYER metal1 ;
  RECT 1768.920 0.000 1770.040 1.120 ;
 END
END A2
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1763.960 0.000 1765.080 1.120 ;
  LAYER metal4 ;
  RECT 1763.960 0.000 1765.080 1.120 ;
  LAYER metal3 ;
  RECT 1763.960 0.000 1765.080 1.120 ;
  LAYER metal2 ;
  RECT 1763.960 0.000 1765.080 1.120 ;
  LAYER metal1 ;
  RECT 1763.960 0.000 1765.080 1.120 ;
 END
END A1
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1761.480 0.000 1762.600 1.120 ;
  LAYER metal4 ;
  RECT 1761.480 0.000 1762.600 1.120 ;
  LAYER metal3 ;
  RECT 1761.480 0.000 1762.600 1.120 ;
  LAYER metal2 ;
  RECT 1761.480 0.000 1762.600 1.120 ;
  LAYER metal1 ;
  RECT 1761.480 0.000 1762.600 1.120 ;
 END
END A0
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1753.420 0.000 1754.540 1.120 ;
  LAYER metal4 ;
  RECT 1753.420 0.000 1754.540 1.120 ;
  LAYER metal3 ;
  RECT 1753.420 0.000 1754.540 1.120 ;
  LAYER metal2 ;
  RECT 1753.420 0.000 1754.540 1.120 ;
  LAYER metal1 ;
  RECT 1753.420 0.000 1754.540 1.120 ;
 END
END A5
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1747.840 0.000 1748.960 1.120 ;
  LAYER metal4 ;
  RECT 1747.840 0.000 1748.960 1.120 ;
  LAYER metal3 ;
  RECT 1747.840 0.000 1748.960 1.120 ;
  LAYER metal2 ;
  RECT 1747.840 0.000 1748.960 1.120 ;
  LAYER metal1 ;
  RECT 1747.840 0.000 1748.960 1.120 ;
 END
END A4
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1741.640 0.000 1742.760 1.120 ;
  LAYER metal4 ;
  RECT 1741.640 0.000 1742.760 1.120 ;
  LAYER metal3 ;
  RECT 1741.640 0.000 1742.760 1.120 ;
  LAYER metal2 ;
  RECT 1741.640 0.000 1742.760 1.120 ;
  LAYER metal1 ;
  RECT 1741.640 0.000 1742.760 1.120 ;
 END
END A3
PIN DIA63
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1719.320 0.000 1720.440 1.120 ;
  LAYER metal4 ;
  RECT 1719.320 0.000 1720.440 1.120 ;
  LAYER metal3 ;
  RECT 1719.320 0.000 1720.440 1.120 ;
  LAYER metal2 ;
  RECT 1719.320 0.000 1720.440 1.120 ;
  LAYER metal1 ;
  RECT 1719.320 0.000 1720.440 1.120 ;
 END
END DIA63
PIN DOA63
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1706.300 0.000 1707.420 1.120 ;
  LAYER metal4 ;
  RECT 1706.300 0.000 1707.420 1.120 ;
  LAYER metal3 ;
  RECT 1706.300 0.000 1707.420 1.120 ;
  LAYER metal2 ;
  RECT 1706.300 0.000 1707.420 1.120 ;
  LAYER metal1 ;
  RECT 1706.300 0.000 1707.420 1.120 ;
 END
END DOA63
PIN DIA62
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1692.660 0.000 1693.780 1.120 ;
  LAYER metal4 ;
  RECT 1692.660 0.000 1693.780 1.120 ;
  LAYER metal3 ;
  RECT 1692.660 0.000 1693.780 1.120 ;
  LAYER metal2 ;
  RECT 1692.660 0.000 1693.780 1.120 ;
  LAYER metal1 ;
  RECT 1692.660 0.000 1693.780 1.120 ;
 END
END DIA62
PIN DOA62
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1679.020 0.000 1680.140 1.120 ;
  LAYER metal4 ;
  RECT 1679.020 0.000 1680.140 1.120 ;
  LAYER metal3 ;
  RECT 1679.020 0.000 1680.140 1.120 ;
  LAYER metal2 ;
  RECT 1679.020 0.000 1680.140 1.120 ;
  LAYER metal1 ;
  RECT 1679.020 0.000 1680.140 1.120 ;
 END
END DOA62
PIN DIA61
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1666.000 0.000 1667.120 1.120 ;
  LAYER metal4 ;
  RECT 1666.000 0.000 1667.120 1.120 ;
  LAYER metal3 ;
  RECT 1666.000 0.000 1667.120 1.120 ;
  LAYER metal2 ;
  RECT 1666.000 0.000 1667.120 1.120 ;
  LAYER metal1 ;
  RECT 1666.000 0.000 1667.120 1.120 ;
 END
END DIA61
PIN DOA61
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1652.360 0.000 1653.480 1.120 ;
  LAYER metal4 ;
  RECT 1652.360 0.000 1653.480 1.120 ;
  LAYER metal3 ;
  RECT 1652.360 0.000 1653.480 1.120 ;
  LAYER metal2 ;
  RECT 1652.360 0.000 1653.480 1.120 ;
  LAYER metal1 ;
  RECT 1652.360 0.000 1653.480 1.120 ;
 END
END DOA61
PIN DIA60
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1638.720 0.000 1639.840 1.120 ;
  LAYER metal4 ;
  RECT 1638.720 0.000 1639.840 1.120 ;
  LAYER metal3 ;
  RECT 1638.720 0.000 1639.840 1.120 ;
  LAYER metal2 ;
  RECT 1638.720 0.000 1639.840 1.120 ;
  LAYER metal1 ;
  RECT 1638.720 0.000 1639.840 1.120 ;
 END
END DIA60
PIN DOA60
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1625.700 0.000 1626.820 1.120 ;
  LAYER metal4 ;
  RECT 1625.700 0.000 1626.820 1.120 ;
  LAYER metal3 ;
  RECT 1625.700 0.000 1626.820 1.120 ;
  LAYER metal2 ;
  RECT 1625.700 0.000 1626.820 1.120 ;
  LAYER metal1 ;
  RECT 1625.700 0.000 1626.820 1.120 ;
 END
END DOA60
PIN DIA59
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1612.060 0.000 1613.180 1.120 ;
  LAYER metal4 ;
  RECT 1612.060 0.000 1613.180 1.120 ;
  LAYER metal3 ;
  RECT 1612.060 0.000 1613.180 1.120 ;
  LAYER metal2 ;
  RECT 1612.060 0.000 1613.180 1.120 ;
  LAYER metal1 ;
  RECT 1612.060 0.000 1613.180 1.120 ;
 END
END DIA59
PIN DOA59
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1598.420 0.000 1599.540 1.120 ;
  LAYER metal4 ;
  RECT 1598.420 0.000 1599.540 1.120 ;
  LAYER metal3 ;
  RECT 1598.420 0.000 1599.540 1.120 ;
  LAYER metal2 ;
  RECT 1598.420 0.000 1599.540 1.120 ;
  LAYER metal1 ;
  RECT 1598.420 0.000 1599.540 1.120 ;
 END
END DOA59
PIN DIA58
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1585.400 0.000 1586.520 1.120 ;
  LAYER metal4 ;
  RECT 1585.400 0.000 1586.520 1.120 ;
  LAYER metal3 ;
  RECT 1585.400 0.000 1586.520 1.120 ;
  LAYER metal2 ;
  RECT 1585.400 0.000 1586.520 1.120 ;
  LAYER metal1 ;
  RECT 1585.400 0.000 1586.520 1.120 ;
 END
END DIA58
PIN DOA58
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1571.760 0.000 1572.880 1.120 ;
  LAYER metal4 ;
  RECT 1571.760 0.000 1572.880 1.120 ;
  LAYER metal3 ;
  RECT 1571.760 0.000 1572.880 1.120 ;
  LAYER metal2 ;
  RECT 1571.760 0.000 1572.880 1.120 ;
  LAYER metal1 ;
  RECT 1571.760 0.000 1572.880 1.120 ;
 END
END DOA58
PIN DIA57
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1558.120 0.000 1559.240 1.120 ;
  LAYER metal4 ;
  RECT 1558.120 0.000 1559.240 1.120 ;
  LAYER metal3 ;
  RECT 1558.120 0.000 1559.240 1.120 ;
  LAYER metal2 ;
  RECT 1558.120 0.000 1559.240 1.120 ;
  LAYER metal1 ;
  RECT 1558.120 0.000 1559.240 1.120 ;
 END
END DIA57
PIN DOA57
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1545.100 0.000 1546.220 1.120 ;
  LAYER metal4 ;
  RECT 1545.100 0.000 1546.220 1.120 ;
  LAYER metal3 ;
  RECT 1545.100 0.000 1546.220 1.120 ;
  LAYER metal2 ;
  RECT 1545.100 0.000 1546.220 1.120 ;
  LAYER metal1 ;
  RECT 1545.100 0.000 1546.220 1.120 ;
 END
END DOA57
PIN DIA56
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1531.460 0.000 1532.580 1.120 ;
  LAYER metal4 ;
  RECT 1531.460 0.000 1532.580 1.120 ;
  LAYER metal3 ;
  RECT 1531.460 0.000 1532.580 1.120 ;
  LAYER metal2 ;
  RECT 1531.460 0.000 1532.580 1.120 ;
  LAYER metal1 ;
  RECT 1531.460 0.000 1532.580 1.120 ;
 END
END DIA56
PIN DOA56
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1517.820 0.000 1518.940 1.120 ;
  LAYER metal4 ;
  RECT 1517.820 0.000 1518.940 1.120 ;
  LAYER metal3 ;
  RECT 1517.820 0.000 1518.940 1.120 ;
  LAYER metal2 ;
  RECT 1517.820 0.000 1518.940 1.120 ;
  LAYER metal1 ;
  RECT 1517.820 0.000 1518.940 1.120 ;
 END
END DOA56
PIN DIA55
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1504.800 0.000 1505.920 1.120 ;
  LAYER metal4 ;
  RECT 1504.800 0.000 1505.920 1.120 ;
  LAYER metal3 ;
  RECT 1504.800 0.000 1505.920 1.120 ;
  LAYER metal2 ;
  RECT 1504.800 0.000 1505.920 1.120 ;
  LAYER metal1 ;
  RECT 1504.800 0.000 1505.920 1.120 ;
 END
END DIA55
PIN DOA55
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1491.160 0.000 1492.280 1.120 ;
  LAYER metal4 ;
  RECT 1491.160 0.000 1492.280 1.120 ;
  LAYER metal3 ;
  RECT 1491.160 0.000 1492.280 1.120 ;
  LAYER metal2 ;
  RECT 1491.160 0.000 1492.280 1.120 ;
  LAYER metal1 ;
  RECT 1491.160 0.000 1492.280 1.120 ;
 END
END DOA55
PIN DIA54
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1477.520 0.000 1478.640 1.120 ;
  LAYER metal4 ;
  RECT 1477.520 0.000 1478.640 1.120 ;
  LAYER metal3 ;
  RECT 1477.520 0.000 1478.640 1.120 ;
  LAYER metal2 ;
  RECT 1477.520 0.000 1478.640 1.120 ;
  LAYER metal1 ;
  RECT 1477.520 0.000 1478.640 1.120 ;
 END
END DIA54
PIN DOA54
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1464.500 0.000 1465.620 1.120 ;
  LAYER metal4 ;
  RECT 1464.500 0.000 1465.620 1.120 ;
  LAYER metal3 ;
  RECT 1464.500 0.000 1465.620 1.120 ;
  LAYER metal2 ;
  RECT 1464.500 0.000 1465.620 1.120 ;
  LAYER metal1 ;
  RECT 1464.500 0.000 1465.620 1.120 ;
 END
END DOA54
PIN DIA53
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1450.860 0.000 1451.980 1.120 ;
  LAYER metal4 ;
  RECT 1450.860 0.000 1451.980 1.120 ;
  LAYER metal3 ;
  RECT 1450.860 0.000 1451.980 1.120 ;
  LAYER metal2 ;
  RECT 1450.860 0.000 1451.980 1.120 ;
  LAYER metal1 ;
  RECT 1450.860 0.000 1451.980 1.120 ;
 END
END DIA53
PIN DOA53
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1437.220 0.000 1438.340 1.120 ;
  LAYER metal4 ;
  RECT 1437.220 0.000 1438.340 1.120 ;
  LAYER metal3 ;
  RECT 1437.220 0.000 1438.340 1.120 ;
  LAYER metal2 ;
  RECT 1437.220 0.000 1438.340 1.120 ;
  LAYER metal1 ;
  RECT 1437.220 0.000 1438.340 1.120 ;
 END
END DOA53
PIN DIA52
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1424.200 0.000 1425.320 1.120 ;
  LAYER metal4 ;
  RECT 1424.200 0.000 1425.320 1.120 ;
  LAYER metal3 ;
  RECT 1424.200 0.000 1425.320 1.120 ;
  LAYER metal2 ;
  RECT 1424.200 0.000 1425.320 1.120 ;
  LAYER metal1 ;
  RECT 1424.200 0.000 1425.320 1.120 ;
 END
END DIA52
PIN DOA52
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1410.560 0.000 1411.680 1.120 ;
  LAYER metal4 ;
  RECT 1410.560 0.000 1411.680 1.120 ;
  LAYER metal3 ;
  RECT 1410.560 0.000 1411.680 1.120 ;
  LAYER metal2 ;
  RECT 1410.560 0.000 1411.680 1.120 ;
  LAYER metal1 ;
  RECT 1410.560 0.000 1411.680 1.120 ;
 END
END DOA52
PIN DIA51
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1396.920 0.000 1398.040 1.120 ;
  LAYER metal4 ;
  RECT 1396.920 0.000 1398.040 1.120 ;
  LAYER metal3 ;
  RECT 1396.920 0.000 1398.040 1.120 ;
  LAYER metal2 ;
  RECT 1396.920 0.000 1398.040 1.120 ;
  LAYER metal1 ;
  RECT 1396.920 0.000 1398.040 1.120 ;
 END
END DIA51
PIN DOA51
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1383.900 0.000 1385.020 1.120 ;
  LAYER metal4 ;
  RECT 1383.900 0.000 1385.020 1.120 ;
  LAYER metal3 ;
  RECT 1383.900 0.000 1385.020 1.120 ;
  LAYER metal2 ;
  RECT 1383.900 0.000 1385.020 1.120 ;
  LAYER metal1 ;
  RECT 1383.900 0.000 1385.020 1.120 ;
 END
END DOA51
PIN DIA50
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1370.260 0.000 1371.380 1.120 ;
  LAYER metal4 ;
  RECT 1370.260 0.000 1371.380 1.120 ;
  LAYER metal3 ;
  RECT 1370.260 0.000 1371.380 1.120 ;
  LAYER metal2 ;
  RECT 1370.260 0.000 1371.380 1.120 ;
  LAYER metal1 ;
  RECT 1370.260 0.000 1371.380 1.120 ;
 END
END DIA50
PIN DOA50
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1356.620 0.000 1357.740 1.120 ;
  LAYER metal4 ;
  RECT 1356.620 0.000 1357.740 1.120 ;
  LAYER metal3 ;
  RECT 1356.620 0.000 1357.740 1.120 ;
  LAYER metal2 ;
  RECT 1356.620 0.000 1357.740 1.120 ;
  LAYER metal1 ;
  RECT 1356.620 0.000 1357.740 1.120 ;
 END
END DOA50
PIN DIA49
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1343.600 0.000 1344.720 1.120 ;
  LAYER metal4 ;
  RECT 1343.600 0.000 1344.720 1.120 ;
  LAYER metal3 ;
  RECT 1343.600 0.000 1344.720 1.120 ;
  LAYER metal2 ;
  RECT 1343.600 0.000 1344.720 1.120 ;
  LAYER metal1 ;
  RECT 1343.600 0.000 1344.720 1.120 ;
 END
END DIA49
PIN DOA49
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1329.960 0.000 1331.080 1.120 ;
  LAYER metal4 ;
  RECT 1329.960 0.000 1331.080 1.120 ;
  LAYER metal3 ;
  RECT 1329.960 0.000 1331.080 1.120 ;
  LAYER metal2 ;
  RECT 1329.960 0.000 1331.080 1.120 ;
  LAYER metal1 ;
  RECT 1329.960 0.000 1331.080 1.120 ;
 END
END DOA49
PIN DIA48
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1316.320 0.000 1317.440 1.120 ;
  LAYER metal4 ;
  RECT 1316.320 0.000 1317.440 1.120 ;
  LAYER metal3 ;
  RECT 1316.320 0.000 1317.440 1.120 ;
  LAYER metal2 ;
  RECT 1316.320 0.000 1317.440 1.120 ;
  LAYER metal1 ;
  RECT 1316.320 0.000 1317.440 1.120 ;
 END
END DIA48
PIN WEAN3
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1305.160 0.000 1306.280 1.120 ;
  LAYER metal4 ;
  RECT 1305.160 0.000 1306.280 1.120 ;
  LAYER metal3 ;
  RECT 1305.160 0.000 1306.280 1.120 ;
  LAYER metal2 ;
  RECT 1305.160 0.000 1306.280 1.120 ;
  LAYER metal1 ;
  RECT 1305.160 0.000 1306.280 1.120 ;
 END
END WEAN3
PIN DOA48
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1302.680 0.000 1303.800 1.120 ;
  LAYER metal4 ;
  RECT 1302.680 0.000 1303.800 1.120 ;
  LAYER metal3 ;
  RECT 1302.680 0.000 1303.800 1.120 ;
  LAYER metal2 ;
  RECT 1302.680 0.000 1303.800 1.120 ;
  LAYER metal1 ;
  RECT 1302.680 0.000 1303.800 1.120 ;
 END
END DOA48
PIN DIA47
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1289.660 0.000 1290.780 1.120 ;
  LAYER metal4 ;
  RECT 1289.660 0.000 1290.780 1.120 ;
  LAYER metal3 ;
  RECT 1289.660 0.000 1290.780 1.120 ;
  LAYER metal2 ;
  RECT 1289.660 0.000 1290.780 1.120 ;
  LAYER metal1 ;
  RECT 1289.660 0.000 1290.780 1.120 ;
 END
END DIA47
PIN DOA47
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1276.020 0.000 1277.140 1.120 ;
  LAYER metal4 ;
  RECT 1276.020 0.000 1277.140 1.120 ;
  LAYER metal3 ;
  RECT 1276.020 0.000 1277.140 1.120 ;
  LAYER metal2 ;
  RECT 1276.020 0.000 1277.140 1.120 ;
  LAYER metal1 ;
  RECT 1276.020 0.000 1277.140 1.120 ;
 END
END DOA47
PIN DIA46
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1262.380 0.000 1263.500 1.120 ;
  LAYER metal4 ;
  RECT 1262.380 0.000 1263.500 1.120 ;
  LAYER metal3 ;
  RECT 1262.380 0.000 1263.500 1.120 ;
  LAYER metal2 ;
  RECT 1262.380 0.000 1263.500 1.120 ;
  LAYER metal1 ;
  RECT 1262.380 0.000 1263.500 1.120 ;
 END
END DIA46
PIN DOA46
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1249.360 0.000 1250.480 1.120 ;
  LAYER metal4 ;
  RECT 1249.360 0.000 1250.480 1.120 ;
  LAYER metal3 ;
  RECT 1249.360 0.000 1250.480 1.120 ;
  LAYER metal2 ;
  RECT 1249.360 0.000 1250.480 1.120 ;
  LAYER metal1 ;
  RECT 1249.360 0.000 1250.480 1.120 ;
 END
END DOA46
PIN DIA45
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1235.720 0.000 1236.840 1.120 ;
  LAYER metal4 ;
  RECT 1235.720 0.000 1236.840 1.120 ;
  LAYER metal3 ;
  RECT 1235.720 0.000 1236.840 1.120 ;
  LAYER metal2 ;
  RECT 1235.720 0.000 1236.840 1.120 ;
  LAYER metal1 ;
  RECT 1235.720 0.000 1236.840 1.120 ;
 END
END DIA45
PIN DOA45
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1222.080 0.000 1223.200 1.120 ;
  LAYER metal4 ;
  RECT 1222.080 0.000 1223.200 1.120 ;
  LAYER metal3 ;
  RECT 1222.080 0.000 1223.200 1.120 ;
  LAYER metal2 ;
  RECT 1222.080 0.000 1223.200 1.120 ;
  LAYER metal1 ;
  RECT 1222.080 0.000 1223.200 1.120 ;
 END
END DOA45
PIN DIA44
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1209.060 0.000 1210.180 1.120 ;
  LAYER metal4 ;
  RECT 1209.060 0.000 1210.180 1.120 ;
  LAYER metal3 ;
  RECT 1209.060 0.000 1210.180 1.120 ;
  LAYER metal2 ;
  RECT 1209.060 0.000 1210.180 1.120 ;
  LAYER metal1 ;
  RECT 1209.060 0.000 1210.180 1.120 ;
 END
END DIA44
PIN DOA44
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1195.420 0.000 1196.540 1.120 ;
  LAYER metal4 ;
  RECT 1195.420 0.000 1196.540 1.120 ;
  LAYER metal3 ;
  RECT 1195.420 0.000 1196.540 1.120 ;
  LAYER metal2 ;
  RECT 1195.420 0.000 1196.540 1.120 ;
  LAYER metal1 ;
  RECT 1195.420 0.000 1196.540 1.120 ;
 END
END DOA44
PIN DIA43
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1181.780 0.000 1182.900 1.120 ;
  LAYER metal4 ;
  RECT 1181.780 0.000 1182.900 1.120 ;
  LAYER metal3 ;
  RECT 1181.780 0.000 1182.900 1.120 ;
  LAYER metal2 ;
  RECT 1181.780 0.000 1182.900 1.120 ;
  LAYER metal1 ;
  RECT 1181.780 0.000 1182.900 1.120 ;
 END
END DIA43
PIN DOA43
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1168.760 0.000 1169.880 1.120 ;
  LAYER metal4 ;
  RECT 1168.760 0.000 1169.880 1.120 ;
  LAYER metal3 ;
  RECT 1168.760 0.000 1169.880 1.120 ;
  LAYER metal2 ;
  RECT 1168.760 0.000 1169.880 1.120 ;
  LAYER metal1 ;
  RECT 1168.760 0.000 1169.880 1.120 ;
 END
END DOA43
PIN DIA42
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1155.120 0.000 1156.240 1.120 ;
  LAYER metal4 ;
  RECT 1155.120 0.000 1156.240 1.120 ;
  LAYER metal3 ;
  RECT 1155.120 0.000 1156.240 1.120 ;
  LAYER metal2 ;
  RECT 1155.120 0.000 1156.240 1.120 ;
  LAYER metal1 ;
  RECT 1155.120 0.000 1156.240 1.120 ;
 END
END DIA42
PIN DOA42
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1141.480 0.000 1142.600 1.120 ;
  LAYER metal4 ;
  RECT 1141.480 0.000 1142.600 1.120 ;
  LAYER metal3 ;
  RECT 1141.480 0.000 1142.600 1.120 ;
  LAYER metal2 ;
  RECT 1141.480 0.000 1142.600 1.120 ;
  LAYER metal1 ;
  RECT 1141.480 0.000 1142.600 1.120 ;
 END
END DOA42
PIN DIA41
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1128.460 0.000 1129.580 1.120 ;
  LAYER metal4 ;
  RECT 1128.460 0.000 1129.580 1.120 ;
  LAYER metal3 ;
  RECT 1128.460 0.000 1129.580 1.120 ;
  LAYER metal2 ;
  RECT 1128.460 0.000 1129.580 1.120 ;
  LAYER metal1 ;
  RECT 1128.460 0.000 1129.580 1.120 ;
 END
END DIA41
PIN DOA41
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1114.820 0.000 1115.940 1.120 ;
  LAYER metal4 ;
  RECT 1114.820 0.000 1115.940 1.120 ;
  LAYER metal3 ;
  RECT 1114.820 0.000 1115.940 1.120 ;
  LAYER metal2 ;
  RECT 1114.820 0.000 1115.940 1.120 ;
  LAYER metal1 ;
  RECT 1114.820 0.000 1115.940 1.120 ;
 END
END DOA41
PIN DIA40
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1101.180 0.000 1102.300 1.120 ;
  LAYER metal4 ;
  RECT 1101.180 0.000 1102.300 1.120 ;
  LAYER metal3 ;
  RECT 1101.180 0.000 1102.300 1.120 ;
  LAYER metal2 ;
  RECT 1101.180 0.000 1102.300 1.120 ;
  LAYER metal1 ;
  RECT 1101.180 0.000 1102.300 1.120 ;
 END
END DIA40
PIN DOA40
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1088.160 0.000 1089.280 1.120 ;
  LAYER metal4 ;
  RECT 1088.160 0.000 1089.280 1.120 ;
  LAYER metal3 ;
  RECT 1088.160 0.000 1089.280 1.120 ;
  LAYER metal2 ;
  RECT 1088.160 0.000 1089.280 1.120 ;
  LAYER metal1 ;
  RECT 1088.160 0.000 1089.280 1.120 ;
 END
END DOA40
PIN DIA39
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1074.520 0.000 1075.640 1.120 ;
  LAYER metal4 ;
  RECT 1074.520 0.000 1075.640 1.120 ;
  LAYER metal3 ;
  RECT 1074.520 0.000 1075.640 1.120 ;
  LAYER metal2 ;
  RECT 1074.520 0.000 1075.640 1.120 ;
  LAYER metal1 ;
  RECT 1074.520 0.000 1075.640 1.120 ;
 END
END DIA39
PIN DOA39
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1060.880 0.000 1062.000 1.120 ;
  LAYER metal4 ;
  RECT 1060.880 0.000 1062.000 1.120 ;
  LAYER metal3 ;
  RECT 1060.880 0.000 1062.000 1.120 ;
  LAYER metal2 ;
  RECT 1060.880 0.000 1062.000 1.120 ;
  LAYER metal1 ;
  RECT 1060.880 0.000 1062.000 1.120 ;
 END
END DOA39
PIN DIA38
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1047.860 0.000 1048.980 1.120 ;
  LAYER metal4 ;
  RECT 1047.860 0.000 1048.980 1.120 ;
  LAYER metal3 ;
  RECT 1047.860 0.000 1048.980 1.120 ;
  LAYER metal2 ;
  RECT 1047.860 0.000 1048.980 1.120 ;
  LAYER metal1 ;
  RECT 1047.860 0.000 1048.980 1.120 ;
 END
END DIA38
PIN DOA38
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1034.220 0.000 1035.340 1.120 ;
  LAYER metal4 ;
  RECT 1034.220 0.000 1035.340 1.120 ;
  LAYER metal3 ;
  RECT 1034.220 0.000 1035.340 1.120 ;
  LAYER metal2 ;
  RECT 1034.220 0.000 1035.340 1.120 ;
  LAYER metal1 ;
  RECT 1034.220 0.000 1035.340 1.120 ;
 END
END DOA38
PIN DIA37
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1020.580 0.000 1021.700 1.120 ;
  LAYER metal4 ;
  RECT 1020.580 0.000 1021.700 1.120 ;
  LAYER metal3 ;
  RECT 1020.580 0.000 1021.700 1.120 ;
  LAYER metal2 ;
  RECT 1020.580 0.000 1021.700 1.120 ;
  LAYER metal1 ;
  RECT 1020.580 0.000 1021.700 1.120 ;
 END
END DIA37
PIN DOA37
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1007.560 0.000 1008.680 1.120 ;
  LAYER metal4 ;
  RECT 1007.560 0.000 1008.680 1.120 ;
  LAYER metal3 ;
  RECT 1007.560 0.000 1008.680 1.120 ;
  LAYER metal2 ;
  RECT 1007.560 0.000 1008.680 1.120 ;
  LAYER metal1 ;
  RECT 1007.560 0.000 1008.680 1.120 ;
 END
END DOA37
PIN DIA36
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 993.920 0.000 995.040 1.120 ;
  LAYER metal4 ;
  RECT 993.920 0.000 995.040 1.120 ;
  LAYER metal3 ;
  RECT 993.920 0.000 995.040 1.120 ;
  LAYER metal2 ;
  RECT 993.920 0.000 995.040 1.120 ;
  LAYER metal1 ;
  RECT 993.920 0.000 995.040 1.120 ;
 END
END DIA36
PIN DOA36
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 980.280 0.000 981.400 1.120 ;
  LAYER metal4 ;
  RECT 980.280 0.000 981.400 1.120 ;
  LAYER metal3 ;
  RECT 980.280 0.000 981.400 1.120 ;
  LAYER metal2 ;
  RECT 980.280 0.000 981.400 1.120 ;
  LAYER metal1 ;
  RECT 980.280 0.000 981.400 1.120 ;
 END
END DOA36
PIN DIA35
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 967.260 0.000 968.380 1.120 ;
  LAYER metal4 ;
  RECT 967.260 0.000 968.380 1.120 ;
  LAYER metal3 ;
  RECT 967.260 0.000 968.380 1.120 ;
  LAYER metal2 ;
  RECT 967.260 0.000 968.380 1.120 ;
  LAYER metal1 ;
  RECT 967.260 0.000 968.380 1.120 ;
 END
END DIA35
PIN DOA35
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 953.620 0.000 954.740 1.120 ;
  LAYER metal4 ;
  RECT 953.620 0.000 954.740 1.120 ;
  LAYER metal3 ;
  RECT 953.620 0.000 954.740 1.120 ;
  LAYER metal2 ;
  RECT 953.620 0.000 954.740 1.120 ;
  LAYER metal1 ;
  RECT 953.620 0.000 954.740 1.120 ;
 END
END DOA35
PIN DIA34
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 939.980 0.000 941.100 1.120 ;
  LAYER metal4 ;
  RECT 939.980 0.000 941.100 1.120 ;
  LAYER metal3 ;
  RECT 939.980 0.000 941.100 1.120 ;
  LAYER metal2 ;
  RECT 939.980 0.000 941.100 1.120 ;
  LAYER metal1 ;
  RECT 939.980 0.000 941.100 1.120 ;
 END
END DIA34
PIN DOA34
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 926.960 0.000 928.080 1.120 ;
  LAYER metal4 ;
  RECT 926.960 0.000 928.080 1.120 ;
  LAYER metal3 ;
  RECT 926.960 0.000 928.080 1.120 ;
  LAYER metal2 ;
  RECT 926.960 0.000 928.080 1.120 ;
  LAYER metal1 ;
  RECT 926.960 0.000 928.080 1.120 ;
 END
END DOA34
PIN DIA33
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 913.320 0.000 914.440 1.120 ;
  LAYER metal4 ;
  RECT 913.320 0.000 914.440 1.120 ;
  LAYER metal3 ;
  RECT 913.320 0.000 914.440 1.120 ;
  LAYER metal2 ;
  RECT 913.320 0.000 914.440 1.120 ;
  LAYER metal1 ;
  RECT 913.320 0.000 914.440 1.120 ;
 END
END DIA33
PIN DOA33
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 899.680 0.000 900.800 1.120 ;
  LAYER metal4 ;
  RECT 899.680 0.000 900.800 1.120 ;
  LAYER metal3 ;
  RECT 899.680 0.000 900.800 1.120 ;
  LAYER metal2 ;
  RECT 899.680 0.000 900.800 1.120 ;
  LAYER metal1 ;
  RECT 899.680 0.000 900.800 1.120 ;
 END
END DOA33
PIN DIA32
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 886.040 0.000 887.160 1.120 ;
  LAYER metal4 ;
  RECT 886.040 0.000 887.160 1.120 ;
  LAYER metal3 ;
  RECT 886.040 0.000 887.160 1.120 ;
  LAYER metal2 ;
  RECT 886.040 0.000 887.160 1.120 ;
  LAYER metal1 ;
  RECT 886.040 0.000 887.160 1.120 ;
 END
END DIA32
PIN WEAN2
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 874.880 0.000 876.000 1.120 ;
  LAYER metal4 ;
  RECT 874.880 0.000 876.000 1.120 ;
  LAYER metal3 ;
  RECT 874.880 0.000 876.000 1.120 ;
  LAYER metal2 ;
  RECT 874.880 0.000 876.000 1.120 ;
  LAYER metal1 ;
  RECT 874.880 0.000 876.000 1.120 ;
 END
END WEAN2
PIN DOA32
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 873.020 0.000 874.140 1.120 ;
  LAYER metal4 ;
  RECT 873.020 0.000 874.140 1.120 ;
  LAYER metal3 ;
  RECT 873.020 0.000 874.140 1.120 ;
  LAYER metal2 ;
  RECT 873.020 0.000 874.140 1.120 ;
  LAYER metal1 ;
  RECT 873.020 0.000 874.140 1.120 ;
 END
END DOA32
PIN DIA31
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 859.380 0.000 860.500 1.120 ;
  LAYER metal4 ;
  RECT 859.380 0.000 860.500 1.120 ;
  LAYER metal3 ;
  RECT 859.380 0.000 860.500 1.120 ;
  LAYER metal2 ;
  RECT 859.380 0.000 860.500 1.120 ;
  LAYER metal1 ;
  RECT 859.380 0.000 860.500 1.120 ;
 END
END DIA31
PIN DOA31
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 845.740 0.000 846.860 1.120 ;
  LAYER metal4 ;
  RECT 845.740 0.000 846.860 1.120 ;
  LAYER metal3 ;
  RECT 845.740 0.000 846.860 1.120 ;
  LAYER metal2 ;
  RECT 845.740 0.000 846.860 1.120 ;
  LAYER metal1 ;
  RECT 845.740 0.000 846.860 1.120 ;
 END
END DOA31
PIN DIA30
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 832.720 0.000 833.840 1.120 ;
  LAYER metal4 ;
  RECT 832.720 0.000 833.840 1.120 ;
  LAYER metal3 ;
  RECT 832.720 0.000 833.840 1.120 ;
  LAYER metal2 ;
  RECT 832.720 0.000 833.840 1.120 ;
  LAYER metal1 ;
  RECT 832.720 0.000 833.840 1.120 ;
 END
END DIA30
PIN DOA30
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 819.080 0.000 820.200 1.120 ;
  LAYER metal4 ;
  RECT 819.080 0.000 820.200 1.120 ;
  LAYER metal3 ;
  RECT 819.080 0.000 820.200 1.120 ;
  LAYER metal2 ;
  RECT 819.080 0.000 820.200 1.120 ;
  LAYER metal1 ;
  RECT 819.080 0.000 820.200 1.120 ;
 END
END DOA30
PIN DIA29
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 805.440 0.000 806.560 1.120 ;
  LAYER metal4 ;
  RECT 805.440 0.000 806.560 1.120 ;
  LAYER metal3 ;
  RECT 805.440 0.000 806.560 1.120 ;
  LAYER metal2 ;
  RECT 805.440 0.000 806.560 1.120 ;
  LAYER metal1 ;
  RECT 805.440 0.000 806.560 1.120 ;
 END
END DIA29
PIN DOA29
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 792.420 0.000 793.540 1.120 ;
  LAYER metal4 ;
  RECT 792.420 0.000 793.540 1.120 ;
  LAYER metal3 ;
  RECT 792.420 0.000 793.540 1.120 ;
  LAYER metal2 ;
  RECT 792.420 0.000 793.540 1.120 ;
  LAYER metal1 ;
  RECT 792.420 0.000 793.540 1.120 ;
 END
END DOA29
PIN DIA28
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 778.780 0.000 779.900 1.120 ;
  LAYER metal4 ;
  RECT 778.780 0.000 779.900 1.120 ;
  LAYER metal3 ;
  RECT 778.780 0.000 779.900 1.120 ;
  LAYER metal2 ;
  RECT 778.780 0.000 779.900 1.120 ;
  LAYER metal1 ;
  RECT 778.780 0.000 779.900 1.120 ;
 END
END DIA28
PIN DOA28
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 765.140 0.000 766.260 1.120 ;
  LAYER metal4 ;
  RECT 765.140 0.000 766.260 1.120 ;
  LAYER metal3 ;
  RECT 765.140 0.000 766.260 1.120 ;
  LAYER metal2 ;
  RECT 765.140 0.000 766.260 1.120 ;
  LAYER metal1 ;
  RECT 765.140 0.000 766.260 1.120 ;
 END
END DOA28
PIN DIA27
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 752.120 0.000 753.240 1.120 ;
  LAYER metal4 ;
  RECT 752.120 0.000 753.240 1.120 ;
  LAYER metal3 ;
  RECT 752.120 0.000 753.240 1.120 ;
  LAYER metal2 ;
  RECT 752.120 0.000 753.240 1.120 ;
  LAYER metal1 ;
  RECT 752.120 0.000 753.240 1.120 ;
 END
END DIA27
PIN DOA27
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 738.480 0.000 739.600 1.120 ;
  LAYER metal4 ;
  RECT 738.480 0.000 739.600 1.120 ;
  LAYER metal3 ;
  RECT 738.480 0.000 739.600 1.120 ;
  LAYER metal2 ;
  RECT 738.480 0.000 739.600 1.120 ;
  LAYER metal1 ;
  RECT 738.480 0.000 739.600 1.120 ;
 END
END DOA27
PIN DIA26
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 724.840 0.000 725.960 1.120 ;
  LAYER metal4 ;
  RECT 724.840 0.000 725.960 1.120 ;
  LAYER metal3 ;
  RECT 724.840 0.000 725.960 1.120 ;
  LAYER metal2 ;
  RECT 724.840 0.000 725.960 1.120 ;
  LAYER metal1 ;
  RECT 724.840 0.000 725.960 1.120 ;
 END
END DIA26
PIN DOA26
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 711.820 0.000 712.940 1.120 ;
  LAYER metal4 ;
  RECT 711.820 0.000 712.940 1.120 ;
  LAYER metal3 ;
  RECT 711.820 0.000 712.940 1.120 ;
  LAYER metal2 ;
  RECT 711.820 0.000 712.940 1.120 ;
  LAYER metal1 ;
  RECT 711.820 0.000 712.940 1.120 ;
 END
END DOA26
PIN DIA25
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 698.180 0.000 699.300 1.120 ;
  LAYER metal4 ;
  RECT 698.180 0.000 699.300 1.120 ;
  LAYER metal3 ;
  RECT 698.180 0.000 699.300 1.120 ;
  LAYER metal2 ;
  RECT 698.180 0.000 699.300 1.120 ;
  LAYER metal1 ;
  RECT 698.180 0.000 699.300 1.120 ;
 END
END DIA25
PIN DOA25
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 684.540 0.000 685.660 1.120 ;
  LAYER metal4 ;
  RECT 684.540 0.000 685.660 1.120 ;
  LAYER metal3 ;
  RECT 684.540 0.000 685.660 1.120 ;
  LAYER metal2 ;
  RECT 684.540 0.000 685.660 1.120 ;
  LAYER metal1 ;
  RECT 684.540 0.000 685.660 1.120 ;
 END
END DOA25
PIN DIA24
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 671.520 0.000 672.640 1.120 ;
  LAYER metal4 ;
  RECT 671.520 0.000 672.640 1.120 ;
  LAYER metal3 ;
  RECT 671.520 0.000 672.640 1.120 ;
  LAYER metal2 ;
  RECT 671.520 0.000 672.640 1.120 ;
  LAYER metal1 ;
  RECT 671.520 0.000 672.640 1.120 ;
 END
END DIA24
PIN DOA24
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 657.880 0.000 659.000 1.120 ;
  LAYER metal4 ;
  RECT 657.880 0.000 659.000 1.120 ;
  LAYER metal3 ;
  RECT 657.880 0.000 659.000 1.120 ;
  LAYER metal2 ;
  RECT 657.880 0.000 659.000 1.120 ;
  LAYER metal1 ;
  RECT 657.880 0.000 659.000 1.120 ;
 END
END DOA24
PIN DIA23
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 644.240 0.000 645.360 1.120 ;
  LAYER metal4 ;
  RECT 644.240 0.000 645.360 1.120 ;
  LAYER metal3 ;
  RECT 644.240 0.000 645.360 1.120 ;
  LAYER metal2 ;
  RECT 644.240 0.000 645.360 1.120 ;
  LAYER metal1 ;
  RECT 644.240 0.000 645.360 1.120 ;
 END
END DIA23
PIN DOA23
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 631.220 0.000 632.340 1.120 ;
  LAYER metal4 ;
  RECT 631.220 0.000 632.340 1.120 ;
  LAYER metal3 ;
  RECT 631.220 0.000 632.340 1.120 ;
  LAYER metal2 ;
  RECT 631.220 0.000 632.340 1.120 ;
  LAYER metal1 ;
  RECT 631.220 0.000 632.340 1.120 ;
 END
END DOA23
PIN DIA22
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 617.580 0.000 618.700 1.120 ;
  LAYER metal4 ;
  RECT 617.580 0.000 618.700 1.120 ;
  LAYER metal3 ;
  RECT 617.580 0.000 618.700 1.120 ;
  LAYER metal2 ;
  RECT 617.580 0.000 618.700 1.120 ;
  LAYER metal1 ;
  RECT 617.580 0.000 618.700 1.120 ;
 END
END DIA22
PIN DOA22
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 603.940 0.000 605.060 1.120 ;
  LAYER metal4 ;
  RECT 603.940 0.000 605.060 1.120 ;
  LAYER metal3 ;
  RECT 603.940 0.000 605.060 1.120 ;
  LAYER metal2 ;
  RECT 603.940 0.000 605.060 1.120 ;
  LAYER metal1 ;
  RECT 603.940 0.000 605.060 1.120 ;
 END
END DOA22
PIN DIA21
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 590.920 0.000 592.040 1.120 ;
  LAYER metal4 ;
  RECT 590.920 0.000 592.040 1.120 ;
  LAYER metal3 ;
  RECT 590.920 0.000 592.040 1.120 ;
  LAYER metal2 ;
  RECT 590.920 0.000 592.040 1.120 ;
  LAYER metal1 ;
  RECT 590.920 0.000 592.040 1.120 ;
 END
END DIA21
PIN DOA21
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 577.280 0.000 578.400 1.120 ;
  LAYER metal4 ;
  RECT 577.280 0.000 578.400 1.120 ;
  LAYER metal3 ;
  RECT 577.280 0.000 578.400 1.120 ;
  LAYER metal2 ;
  RECT 577.280 0.000 578.400 1.120 ;
  LAYER metal1 ;
  RECT 577.280 0.000 578.400 1.120 ;
 END
END DOA21
PIN DIA20
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 563.640 0.000 564.760 1.120 ;
  LAYER metal4 ;
  RECT 563.640 0.000 564.760 1.120 ;
  LAYER metal3 ;
  RECT 563.640 0.000 564.760 1.120 ;
  LAYER metal2 ;
  RECT 563.640 0.000 564.760 1.120 ;
  LAYER metal1 ;
  RECT 563.640 0.000 564.760 1.120 ;
 END
END DIA20
PIN DOA20
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 550.620 0.000 551.740 1.120 ;
  LAYER metal4 ;
  RECT 550.620 0.000 551.740 1.120 ;
  LAYER metal3 ;
  RECT 550.620 0.000 551.740 1.120 ;
  LAYER metal2 ;
  RECT 550.620 0.000 551.740 1.120 ;
  LAYER metal1 ;
  RECT 550.620 0.000 551.740 1.120 ;
 END
END DOA20
PIN DIA19
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 536.980 0.000 538.100 1.120 ;
  LAYER metal4 ;
  RECT 536.980 0.000 538.100 1.120 ;
  LAYER metal3 ;
  RECT 536.980 0.000 538.100 1.120 ;
  LAYER metal2 ;
  RECT 536.980 0.000 538.100 1.120 ;
  LAYER metal1 ;
  RECT 536.980 0.000 538.100 1.120 ;
 END
END DIA19
PIN DOA19
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 523.340 0.000 524.460 1.120 ;
  LAYER metal4 ;
  RECT 523.340 0.000 524.460 1.120 ;
  LAYER metal3 ;
  RECT 523.340 0.000 524.460 1.120 ;
  LAYER metal2 ;
  RECT 523.340 0.000 524.460 1.120 ;
  LAYER metal1 ;
  RECT 523.340 0.000 524.460 1.120 ;
 END
END DOA19
PIN DIA18
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 510.320 0.000 511.440 1.120 ;
  LAYER metal4 ;
  RECT 510.320 0.000 511.440 1.120 ;
  LAYER metal3 ;
  RECT 510.320 0.000 511.440 1.120 ;
  LAYER metal2 ;
  RECT 510.320 0.000 511.440 1.120 ;
  LAYER metal1 ;
  RECT 510.320 0.000 511.440 1.120 ;
 END
END DIA18
PIN DOA18
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 496.680 0.000 497.800 1.120 ;
  LAYER metal4 ;
  RECT 496.680 0.000 497.800 1.120 ;
  LAYER metal3 ;
  RECT 496.680 0.000 497.800 1.120 ;
  LAYER metal2 ;
  RECT 496.680 0.000 497.800 1.120 ;
  LAYER metal1 ;
  RECT 496.680 0.000 497.800 1.120 ;
 END
END DOA18
PIN DIA17
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 483.040 0.000 484.160 1.120 ;
  LAYER metal4 ;
  RECT 483.040 0.000 484.160 1.120 ;
  LAYER metal3 ;
  RECT 483.040 0.000 484.160 1.120 ;
  LAYER metal2 ;
  RECT 483.040 0.000 484.160 1.120 ;
  LAYER metal1 ;
  RECT 483.040 0.000 484.160 1.120 ;
 END
END DIA17
PIN DOA17
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 469.400 0.000 470.520 1.120 ;
  LAYER metal4 ;
  RECT 469.400 0.000 470.520 1.120 ;
  LAYER metal3 ;
  RECT 469.400 0.000 470.520 1.120 ;
  LAYER metal2 ;
  RECT 469.400 0.000 470.520 1.120 ;
  LAYER metal1 ;
  RECT 469.400 0.000 470.520 1.120 ;
 END
END DOA17
PIN DIA16
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 456.380 0.000 457.500 1.120 ;
  LAYER metal4 ;
  RECT 456.380 0.000 457.500 1.120 ;
  LAYER metal3 ;
  RECT 456.380 0.000 457.500 1.120 ;
  LAYER metal2 ;
  RECT 456.380 0.000 457.500 1.120 ;
  LAYER metal1 ;
  RECT 456.380 0.000 457.500 1.120 ;
 END
END DIA16
PIN WEAN1
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 445.220 0.000 446.340 1.120 ;
  LAYER metal4 ;
  RECT 445.220 0.000 446.340 1.120 ;
  LAYER metal3 ;
  RECT 445.220 0.000 446.340 1.120 ;
  LAYER metal2 ;
  RECT 445.220 0.000 446.340 1.120 ;
  LAYER metal1 ;
  RECT 445.220 0.000 446.340 1.120 ;
 END
END WEAN1
PIN DOA16
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 442.740 0.000 443.860 1.120 ;
  LAYER metal4 ;
  RECT 442.740 0.000 443.860 1.120 ;
  LAYER metal3 ;
  RECT 442.740 0.000 443.860 1.120 ;
  LAYER metal2 ;
  RECT 442.740 0.000 443.860 1.120 ;
  LAYER metal1 ;
  RECT 442.740 0.000 443.860 1.120 ;
 END
END DOA16
PIN DIA15
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER metal4 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER metal3 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER metal2 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER metal1 ;
  RECT 429.100 0.000 430.220 1.120 ;
 END
END DIA15
PIN DOA15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 416.080 0.000 417.200 1.120 ;
  LAYER metal4 ;
  RECT 416.080 0.000 417.200 1.120 ;
  LAYER metal3 ;
  RECT 416.080 0.000 417.200 1.120 ;
  LAYER metal2 ;
  RECT 416.080 0.000 417.200 1.120 ;
  LAYER metal1 ;
  RECT 416.080 0.000 417.200 1.120 ;
 END
END DOA15
PIN DIA14
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER metal4 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER metal3 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER metal2 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER metal1 ;
  RECT 402.440 0.000 403.560 1.120 ;
 END
END DIA14
PIN DOA14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 388.800 0.000 389.920 1.120 ;
  LAYER metal4 ;
  RECT 388.800 0.000 389.920 1.120 ;
  LAYER metal3 ;
  RECT 388.800 0.000 389.920 1.120 ;
  LAYER metal2 ;
  RECT 388.800 0.000 389.920 1.120 ;
  LAYER metal1 ;
  RECT 388.800 0.000 389.920 1.120 ;
 END
END DOA14
PIN DIA13
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 375.780 0.000 376.900 1.120 ;
  LAYER metal4 ;
  RECT 375.780 0.000 376.900 1.120 ;
  LAYER metal3 ;
  RECT 375.780 0.000 376.900 1.120 ;
  LAYER metal2 ;
  RECT 375.780 0.000 376.900 1.120 ;
  LAYER metal1 ;
  RECT 375.780 0.000 376.900 1.120 ;
 END
END DIA13
PIN DOA13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 362.140 0.000 363.260 1.120 ;
  LAYER metal4 ;
  RECT 362.140 0.000 363.260 1.120 ;
  LAYER metal3 ;
  RECT 362.140 0.000 363.260 1.120 ;
  LAYER metal2 ;
  RECT 362.140 0.000 363.260 1.120 ;
  LAYER metal1 ;
  RECT 362.140 0.000 363.260 1.120 ;
 END
END DOA13
PIN DIA12
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER metal4 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER metal3 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER metal2 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER metal1 ;
  RECT 348.500 0.000 349.620 1.120 ;
 END
END DIA12
PIN DOA12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 335.480 0.000 336.600 1.120 ;
  LAYER metal4 ;
  RECT 335.480 0.000 336.600 1.120 ;
  LAYER metal3 ;
  RECT 335.480 0.000 336.600 1.120 ;
  LAYER metal2 ;
  RECT 335.480 0.000 336.600 1.120 ;
  LAYER metal1 ;
  RECT 335.480 0.000 336.600 1.120 ;
 END
END DOA12
PIN DIA11
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 321.840 0.000 322.960 1.120 ;
  LAYER metal4 ;
  RECT 321.840 0.000 322.960 1.120 ;
  LAYER metal3 ;
  RECT 321.840 0.000 322.960 1.120 ;
  LAYER metal2 ;
  RECT 321.840 0.000 322.960 1.120 ;
  LAYER metal1 ;
  RECT 321.840 0.000 322.960 1.120 ;
 END
END DIA11
PIN DOA11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 308.200 0.000 309.320 1.120 ;
  LAYER metal4 ;
  RECT 308.200 0.000 309.320 1.120 ;
  LAYER metal3 ;
  RECT 308.200 0.000 309.320 1.120 ;
  LAYER metal2 ;
  RECT 308.200 0.000 309.320 1.120 ;
  LAYER metal1 ;
  RECT 308.200 0.000 309.320 1.120 ;
 END
END DOA11
PIN DIA10
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 295.180 0.000 296.300 1.120 ;
  LAYER metal4 ;
  RECT 295.180 0.000 296.300 1.120 ;
  LAYER metal3 ;
  RECT 295.180 0.000 296.300 1.120 ;
  LAYER metal2 ;
  RECT 295.180 0.000 296.300 1.120 ;
  LAYER metal1 ;
  RECT 295.180 0.000 296.300 1.120 ;
 END
END DIA10
PIN DOA10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 281.540 0.000 282.660 1.120 ;
  LAYER metal4 ;
  RECT 281.540 0.000 282.660 1.120 ;
  LAYER metal3 ;
  RECT 281.540 0.000 282.660 1.120 ;
  LAYER metal2 ;
  RECT 281.540 0.000 282.660 1.120 ;
  LAYER metal1 ;
  RECT 281.540 0.000 282.660 1.120 ;
 END
END DOA10
PIN DIA9
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal4 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal3 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal2 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal1 ;
  RECT 267.900 0.000 269.020 1.120 ;
 END
END DIA9
PIN DOA9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER metal4 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER metal3 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER metal2 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER metal1 ;
  RECT 254.880 0.000 256.000 1.120 ;
 END
END DOA9
PIN DIA8
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal4 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal3 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal2 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal1 ;
  RECT 241.240 0.000 242.360 1.120 ;
 END
END DIA8
PIN DOA8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 227.600 0.000 228.720 1.120 ;
  LAYER metal4 ;
  RECT 227.600 0.000 228.720 1.120 ;
  LAYER metal3 ;
  RECT 227.600 0.000 228.720 1.120 ;
  LAYER metal2 ;
  RECT 227.600 0.000 228.720 1.120 ;
  LAYER metal1 ;
  RECT 227.600 0.000 228.720 1.120 ;
 END
END DOA8
PIN DIA7
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 214.580 0.000 215.700 1.120 ;
  LAYER metal4 ;
  RECT 214.580 0.000 215.700 1.120 ;
  LAYER metal3 ;
  RECT 214.580 0.000 215.700 1.120 ;
  LAYER metal2 ;
  RECT 214.580 0.000 215.700 1.120 ;
  LAYER metal1 ;
  RECT 214.580 0.000 215.700 1.120 ;
 END
END DIA7
PIN DOA7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 200.940 0.000 202.060 1.120 ;
  LAYER metal4 ;
  RECT 200.940 0.000 202.060 1.120 ;
  LAYER metal3 ;
  RECT 200.940 0.000 202.060 1.120 ;
  LAYER metal2 ;
  RECT 200.940 0.000 202.060 1.120 ;
  LAYER metal1 ;
  RECT 200.940 0.000 202.060 1.120 ;
 END
END DOA7
PIN DIA6
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER metal4 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER metal3 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER metal2 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER metal1 ;
  RECT 187.300 0.000 188.420 1.120 ;
 END
END DIA6
PIN DOA6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 174.280 0.000 175.400 1.120 ;
  LAYER metal4 ;
  RECT 174.280 0.000 175.400 1.120 ;
  LAYER metal3 ;
  RECT 174.280 0.000 175.400 1.120 ;
  LAYER metal2 ;
  RECT 174.280 0.000 175.400 1.120 ;
  LAYER metal1 ;
  RECT 174.280 0.000 175.400 1.120 ;
 END
END DOA6
PIN DIA5
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 160.640 0.000 161.760 1.120 ;
  LAYER metal4 ;
  RECT 160.640 0.000 161.760 1.120 ;
  LAYER metal3 ;
  RECT 160.640 0.000 161.760 1.120 ;
  LAYER metal2 ;
  RECT 160.640 0.000 161.760 1.120 ;
  LAYER metal1 ;
  RECT 160.640 0.000 161.760 1.120 ;
 END
END DIA5
PIN DOA5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 147.000 0.000 148.120 1.120 ;
  LAYER metal4 ;
  RECT 147.000 0.000 148.120 1.120 ;
  LAYER metal3 ;
  RECT 147.000 0.000 148.120 1.120 ;
  LAYER metal2 ;
  RECT 147.000 0.000 148.120 1.120 ;
  LAYER metal1 ;
  RECT 147.000 0.000 148.120 1.120 ;
 END
END DOA5
PIN DIA4
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER metal4 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER metal3 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER metal2 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER metal1 ;
  RECT 133.980 0.000 135.100 1.120 ;
 END
END DIA4
PIN DOA4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 120.340 0.000 121.460 1.120 ;
  LAYER metal4 ;
  RECT 120.340 0.000 121.460 1.120 ;
  LAYER metal3 ;
  RECT 120.340 0.000 121.460 1.120 ;
  LAYER metal2 ;
  RECT 120.340 0.000 121.460 1.120 ;
  LAYER metal1 ;
  RECT 120.340 0.000 121.460 1.120 ;
 END
END DOA4
PIN DIA3
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal4 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal3 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal2 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal1 ;
  RECT 106.700 0.000 107.820 1.120 ;
 END
END DIA3
PIN DOA3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 93.680 0.000 94.800 1.120 ;
  LAYER metal4 ;
  RECT 93.680 0.000 94.800 1.120 ;
  LAYER metal3 ;
  RECT 93.680 0.000 94.800 1.120 ;
  LAYER metal2 ;
  RECT 93.680 0.000 94.800 1.120 ;
  LAYER metal1 ;
  RECT 93.680 0.000 94.800 1.120 ;
 END
END DOA3
PIN DIA2
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 80.040 0.000 81.160 1.120 ;
  LAYER metal4 ;
  RECT 80.040 0.000 81.160 1.120 ;
  LAYER metal3 ;
  RECT 80.040 0.000 81.160 1.120 ;
  LAYER metal2 ;
  RECT 80.040 0.000 81.160 1.120 ;
  LAYER metal1 ;
  RECT 80.040 0.000 81.160 1.120 ;
 END
END DIA2
PIN DOA2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 66.400 0.000 67.520 1.120 ;
  LAYER metal4 ;
  RECT 66.400 0.000 67.520 1.120 ;
  LAYER metal3 ;
  RECT 66.400 0.000 67.520 1.120 ;
  LAYER metal2 ;
  RECT 66.400 0.000 67.520 1.120 ;
  LAYER metal1 ;
  RECT 66.400 0.000 67.520 1.120 ;
 END
END DOA2
PIN DIA1
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER metal4 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER metal3 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER metal2 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER metal1 ;
  RECT 52.760 0.000 53.880 1.120 ;
 END
END DIA1
PIN DOA1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER metal4 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER metal3 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER metal2 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER metal1 ;
  RECT 39.740 0.000 40.860 1.120 ;
 END
END DOA1
PIN DIA0
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER metal4 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER metal3 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER metal2 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER metal1 ;
  RECT 26.100 0.000 27.220 1.120 ;
 END
END DIA0
PIN WEAN0
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 14.940 0.000 16.060 1.120 ;
  LAYER metal4 ;
  RECT 14.940 0.000 16.060 1.120 ;
  LAYER metal3 ;
  RECT 14.940 0.000 16.060 1.120 ;
  LAYER metal2 ;
  RECT 14.940 0.000 16.060 1.120 ;
  LAYER metal1 ;
  RECT 14.940 0.000 16.060 1.120 ;
 END
END WEAN0
PIN DOA0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER metal4 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER metal3 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER metal2 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER metal1 ;
  RECT 12.460 0.000 13.580 1.120 ;
 END
END DOA0
OBS
  LAYER metal1 SPACING 0.280 ;
  RECT 0.000 0.140 3547.640 179.620 ;
  LAYER metal2 SPACING 0.320 ;
  RECT 0.000 0.140 3547.640 179.620 ;
  LAYER metal3 SPACING 0.320 ;
  RECT 0.000 0.140 3547.640 179.620 ;
  LAYER metal4 SPACING 0.600 ;
  RECT 0.000 0.140 3547.640 179.620 ;
  LAYER via ;
  RECT 0.000 0.140 3547.640 179.620 ;
  LAYER via2 ;
  RECT 0.000 0.140 3547.640 179.620 ;
  LAYER via3 ;
  RECT 0.000 0.140 3547.640 179.620 ;
END
END word64
END LIBRARY



