`timescale 1ns/10ps
module cnn_top(
	clk,
	rst,
	input_data,
	predict_result
);
