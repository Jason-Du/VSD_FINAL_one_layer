`ifndef DEF_SVH
`define DEF_SVH

`define WORDLENGTH 16
`define LAYER1_WIDTH 32
`define LAYER1_SET_COUNT `LAYER1_WIDTH*2+3-1
`define LAYER1_OUTPUT_LENGTH 128
`define LAYER1_WEIGHT_INPUT_LENGTH 48
`define LAYER1_OUTPUT_CHANNEL_NUM 8
`define LAYER1_SYSTOLIC_WEIGHT_NUM `LAYER1_OUTPUT_CHANNEL_NUM*9

`define LAYER2_WIDTH 30
`define LAYER2_SET_COUNT `LAYER2_WIDTH*2+3-1 
`define LAYER2_OUTPUT_LENGTH 128
`define LAYER2_WEIGHT_INPUT_LENGTH 128
`define LAYER2_OUTPUT_CHANNEL_NUM 8
`define LAYER2_SYSTOLIC_WEIGHT_NUM `LAYER1_OUTPUT_CHANNEL_NUM*9


`define LAYER3_WIDTH 28
`define LAYER3_SET_COUNT `LAYER3_WIDTH*1+2-1 
`define LAYER3_OUTPUT_LENGTH 128

`define LAYER3_WEIGHT_INPUT_LENGTH 128
/*
`define LAYER3_OUTPUT_CHANNEL_NUM 8
`define LAYER3_SYSTOLIC_WEIGHT_NUM `LAYER1_OUTPUT_CHANNEL_NUM*9
*/


`endif