module counter(



);