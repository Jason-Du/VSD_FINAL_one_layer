# 
#              Synchronous Dual Port SRAM Compiler 
# 
#                    UMC 0.18um Generic Logic Process 
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : pixel_sram
#       Words            : 1024
#       Bits             : 16
#       Byte-Write       : 3
#       Aspect Ratio     : 1
#       Output Loading   : 0.5  (pf)
#       Data Slew        : 0.5  (ns)
#       CK Slew          : 0.5  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2021/01/06 16:25:19
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO pixel_sram
CLASS BLOCK ;
FOREIGN pixel_sram 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 1445.840 BY 544.320 ;
SYMMETRY x y r90 ;
SITE core ;
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal5 ;
  RECT 1444.720 521.140 1445.840 524.380 ;
  LAYER metal4 ;
  RECT 1444.720 521.140 1445.840 524.380 ;
  LAYER metal3 ;
  RECT 1444.720 521.140 1445.840 524.380 ;
  LAYER metal2 ;
  RECT 1444.720 521.140 1445.840 524.380 ;
  LAYER metal1 ;
  RECT 1444.720 521.140 1445.840 524.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 513.300 1445.840 516.540 ;
  LAYER metal4 ;
  RECT 1444.720 513.300 1445.840 516.540 ;
  LAYER metal3 ;
  RECT 1444.720 513.300 1445.840 516.540 ;
  LAYER metal2 ;
  RECT 1444.720 513.300 1445.840 516.540 ;
  LAYER metal1 ;
  RECT 1444.720 513.300 1445.840 516.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 505.460 1445.840 508.700 ;
  LAYER metal4 ;
  RECT 1444.720 505.460 1445.840 508.700 ;
  LAYER metal3 ;
  RECT 1444.720 505.460 1445.840 508.700 ;
  LAYER metal2 ;
  RECT 1444.720 505.460 1445.840 508.700 ;
  LAYER metal1 ;
  RECT 1444.720 505.460 1445.840 508.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 497.620 1445.840 500.860 ;
  LAYER metal4 ;
  RECT 1444.720 497.620 1445.840 500.860 ;
  LAYER metal3 ;
  RECT 1444.720 497.620 1445.840 500.860 ;
  LAYER metal2 ;
  RECT 1444.720 497.620 1445.840 500.860 ;
  LAYER metal1 ;
  RECT 1444.720 497.620 1445.840 500.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 489.780 1445.840 493.020 ;
  LAYER metal4 ;
  RECT 1444.720 489.780 1445.840 493.020 ;
  LAYER metal3 ;
  RECT 1444.720 489.780 1445.840 493.020 ;
  LAYER metal2 ;
  RECT 1444.720 489.780 1445.840 493.020 ;
  LAYER metal1 ;
  RECT 1444.720 489.780 1445.840 493.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 481.940 1445.840 485.180 ;
  LAYER metal4 ;
  RECT 1444.720 481.940 1445.840 485.180 ;
  LAYER metal3 ;
  RECT 1444.720 481.940 1445.840 485.180 ;
  LAYER metal2 ;
  RECT 1444.720 481.940 1445.840 485.180 ;
  LAYER metal1 ;
  RECT 1444.720 481.940 1445.840 485.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 442.740 1445.840 445.980 ;
  LAYER metal4 ;
  RECT 1444.720 442.740 1445.840 445.980 ;
  LAYER metal3 ;
  RECT 1444.720 442.740 1445.840 445.980 ;
  LAYER metal2 ;
  RECT 1444.720 442.740 1445.840 445.980 ;
  LAYER metal1 ;
  RECT 1444.720 442.740 1445.840 445.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 434.900 1445.840 438.140 ;
  LAYER metal4 ;
  RECT 1444.720 434.900 1445.840 438.140 ;
  LAYER metal3 ;
  RECT 1444.720 434.900 1445.840 438.140 ;
  LAYER metal2 ;
  RECT 1444.720 434.900 1445.840 438.140 ;
  LAYER metal1 ;
  RECT 1444.720 434.900 1445.840 438.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 427.060 1445.840 430.300 ;
  LAYER metal4 ;
  RECT 1444.720 427.060 1445.840 430.300 ;
  LAYER metal3 ;
  RECT 1444.720 427.060 1445.840 430.300 ;
  LAYER metal2 ;
  RECT 1444.720 427.060 1445.840 430.300 ;
  LAYER metal1 ;
  RECT 1444.720 427.060 1445.840 430.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 419.220 1445.840 422.460 ;
  LAYER metal4 ;
  RECT 1444.720 419.220 1445.840 422.460 ;
  LAYER metal3 ;
  RECT 1444.720 419.220 1445.840 422.460 ;
  LAYER metal2 ;
  RECT 1444.720 419.220 1445.840 422.460 ;
  LAYER metal1 ;
  RECT 1444.720 419.220 1445.840 422.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 411.380 1445.840 414.620 ;
  LAYER metal4 ;
  RECT 1444.720 411.380 1445.840 414.620 ;
  LAYER metal3 ;
  RECT 1444.720 411.380 1445.840 414.620 ;
  LAYER metal2 ;
  RECT 1444.720 411.380 1445.840 414.620 ;
  LAYER metal1 ;
  RECT 1444.720 411.380 1445.840 414.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 403.540 1445.840 406.780 ;
  LAYER metal4 ;
  RECT 1444.720 403.540 1445.840 406.780 ;
  LAYER metal3 ;
  RECT 1444.720 403.540 1445.840 406.780 ;
  LAYER metal2 ;
  RECT 1444.720 403.540 1445.840 406.780 ;
  LAYER metal1 ;
  RECT 1444.720 403.540 1445.840 406.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 364.340 1445.840 367.580 ;
  LAYER metal4 ;
  RECT 1444.720 364.340 1445.840 367.580 ;
  LAYER metal3 ;
  RECT 1444.720 364.340 1445.840 367.580 ;
  LAYER metal2 ;
  RECT 1444.720 364.340 1445.840 367.580 ;
  LAYER metal1 ;
  RECT 1444.720 364.340 1445.840 367.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 356.500 1445.840 359.740 ;
  LAYER metal4 ;
  RECT 1444.720 356.500 1445.840 359.740 ;
  LAYER metal3 ;
  RECT 1444.720 356.500 1445.840 359.740 ;
  LAYER metal2 ;
  RECT 1444.720 356.500 1445.840 359.740 ;
  LAYER metal1 ;
  RECT 1444.720 356.500 1445.840 359.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 348.660 1445.840 351.900 ;
  LAYER metal4 ;
  RECT 1444.720 348.660 1445.840 351.900 ;
  LAYER metal3 ;
  RECT 1444.720 348.660 1445.840 351.900 ;
  LAYER metal2 ;
  RECT 1444.720 348.660 1445.840 351.900 ;
  LAYER metal1 ;
  RECT 1444.720 348.660 1445.840 351.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 340.820 1445.840 344.060 ;
  LAYER metal4 ;
  RECT 1444.720 340.820 1445.840 344.060 ;
  LAYER metal3 ;
  RECT 1444.720 340.820 1445.840 344.060 ;
  LAYER metal2 ;
  RECT 1444.720 340.820 1445.840 344.060 ;
  LAYER metal1 ;
  RECT 1444.720 340.820 1445.840 344.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 332.980 1445.840 336.220 ;
  LAYER metal4 ;
  RECT 1444.720 332.980 1445.840 336.220 ;
  LAYER metal3 ;
  RECT 1444.720 332.980 1445.840 336.220 ;
  LAYER metal2 ;
  RECT 1444.720 332.980 1445.840 336.220 ;
  LAYER metal1 ;
  RECT 1444.720 332.980 1445.840 336.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 325.140 1445.840 328.380 ;
  LAYER metal4 ;
  RECT 1444.720 325.140 1445.840 328.380 ;
  LAYER metal3 ;
  RECT 1444.720 325.140 1445.840 328.380 ;
  LAYER metal2 ;
  RECT 1444.720 325.140 1445.840 328.380 ;
  LAYER metal1 ;
  RECT 1444.720 325.140 1445.840 328.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 285.940 1445.840 289.180 ;
  LAYER metal4 ;
  RECT 1444.720 285.940 1445.840 289.180 ;
  LAYER metal3 ;
  RECT 1444.720 285.940 1445.840 289.180 ;
  LAYER metal2 ;
  RECT 1444.720 285.940 1445.840 289.180 ;
  LAYER metal1 ;
  RECT 1444.720 285.940 1445.840 289.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 278.100 1445.840 281.340 ;
  LAYER metal4 ;
  RECT 1444.720 278.100 1445.840 281.340 ;
  LAYER metal3 ;
  RECT 1444.720 278.100 1445.840 281.340 ;
  LAYER metal2 ;
  RECT 1444.720 278.100 1445.840 281.340 ;
  LAYER metal1 ;
  RECT 1444.720 278.100 1445.840 281.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 270.260 1445.840 273.500 ;
  LAYER metal4 ;
  RECT 1444.720 270.260 1445.840 273.500 ;
  LAYER metal3 ;
  RECT 1444.720 270.260 1445.840 273.500 ;
  LAYER metal2 ;
  RECT 1444.720 270.260 1445.840 273.500 ;
  LAYER metal1 ;
  RECT 1444.720 270.260 1445.840 273.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 262.420 1445.840 265.660 ;
  LAYER metal4 ;
  RECT 1444.720 262.420 1445.840 265.660 ;
  LAYER metal3 ;
  RECT 1444.720 262.420 1445.840 265.660 ;
  LAYER metal2 ;
  RECT 1444.720 262.420 1445.840 265.660 ;
  LAYER metal1 ;
  RECT 1444.720 262.420 1445.840 265.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 254.580 1445.840 257.820 ;
  LAYER metal4 ;
  RECT 1444.720 254.580 1445.840 257.820 ;
  LAYER metal3 ;
  RECT 1444.720 254.580 1445.840 257.820 ;
  LAYER metal2 ;
  RECT 1444.720 254.580 1445.840 257.820 ;
  LAYER metal1 ;
  RECT 1444.720 254.580 1445.840 257.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 246.740 1445.840 249.980 ;
  LAYER metal4 ;
  RECT 1444.720 246.740 1445.840 249.980 ;
  LAYER metal3 ;
  RECT 1444.720 246.740 1445.840 249.980 ;
  LAYER metal2 ;
  RECT 1444.720 246.740 1445.840 249.980 ;
  LAYER metal1 ;
  RECT 1444.720 246.740 1445.840 249.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 207.540 1445.840 210.780 ;
  LAYER metal4 ;
  RECT 1444.720 207.540 1445.840 210.780 ;
  LAYER metal3 ;
  RECT 1444.720 207.540 1445.840 210.780 ;
  LAYER metal2 ;
  RECT 1444.720 207.540 1445.840 210.780 ;
  LAYER metal1 ;
  RECT 1444.720 207.540 1445.840 210.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 199.700 1445.840 202.940 ;
  LAYER metal4 ;
  RECT 1444.720 199.700 1445.840 202.940 ;
  LAYER metal3 ;
  RECT 1444.720 199.700 1445.840 202.940 ;
  LAYER metal2 ;
  RECT 1444.720 199.700 1445.840 202.940 ;
  LAYER metal1 ;
  RECT 1444.720 199.700 1445.840 202.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 191.860 1445.840 195.100 ;
  LAYER metal4 ;
  RECT 1444.720 191.860 1445.840 195.100 ;
  LAYER metal3 ;
  RECT 1444.720 191.860 1445.840 195.100 ;
  LAYER metal2 ;
  RECT 1444.720 191.860 1445.840 195.100 ;
  LAYER metal1 ;
  RECT 1444.720 191.860 1445.840 195.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 184.020 1445.840 187.260 ;
  LAYER metal4 ;
  RECT 1444.720 184.020 1445.840 187.260 ;
  LAYER metal3 ;
  RECT 1444.720 184.020 1445.840 187.260 ;
  LAYER metal2 ;
  RECT 1444.720 184.020 1445.840 187.260 ;
  LAYER metal1 ;
  RECT 1444.720 184.020 1445.840 187.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 176.180 1445.840 179.420 ;
  LAYER metal4 ;
  RECT 1444.720 176.180 1445.840 179.420 ;
  LAYER metal3 ;
  RECT 1444.720 176.180 1445.840 179.420 ;
  LAYER metal2 ;
  RECT 1444.720 176.180 1445.840 179.420 ;
  LAYER metal1 ;
  RECT 1444.720 176.180 1445.840 179.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 168.340 1445.840 171.580 ;
  LAYER metal4 ;
  RECT 1444.720 168.340 1445.840 171.580 ;
  LAYER metal3 ;
  RECT 1444.720 168.340 1445.840 171.580 ;
  LAYER metal2 ;
  RECT 1444.720 168.340 1445.840 171.580 ;
  LAYER metal1 ;
  RECT 1444.720 168.340 1445.840 171.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 129.140 1445.840 132.380 ;
  LAYER metal4 ;
  RECT 1444.720 129.140 1445.840 132.380 ;
  LAYER metal3 ;
  RECT 1444.720 129.140 1445.840 132.380 ;
  LAYER metal2 ;
  RECT 1444.720 129.140 1445.840 132.380 ;
  LAYER metal1 ;
  RECT 1444.720 129.140 1445.840 132.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 121.300 1445.840 124.540 ;
  LAYER metal4 ;
  RECT 1444.720 121.300 1445.840 124.540 ;
  LAYER metal3 ;
  RECT 1444.720 121.300 1445.840 124.540 ;
  LAYER metal2 ;
  RECT 1444.720 121.300 1445.840 124.540 ;
  LAYER metal1 ;
  RECT 1444.720 121.300 1445.840 124.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 113.460 1445.840 116.700 ;
  LAYER metal4 ;
  RECT 1444.720 113.460 1445.840 116.700 ;
  LAYER metal3 ;
  RECT 1444.720 113.460 1445.840 116.700 ;
  LAYER metal2 ;
  RECT 1444.720 113.460 1445.840 116.700 ;
  LAYER metal1 ;
  RECT 1444.720 113.460 1445.840 116.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 105.620 1445.840 108.860 ;
  LAYER metal4 ;
  RECT 1444.720 105.620 1445.840 108.860 ;
  LAYER metal3 ;
  RECT 1444.720 105.620 1445.840 108.860 ;
  LAYER metal2 ;
  RECT 1444.720 105.620 1445.840 108.860 ;
  LAYER metal1 ;
  RECT 1444.720 105.620 1445.840 108.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 97.780 1445.840 101.020 ;
  LAYER metal4 ;
  RECT 1444.720 97.780 1445.840 101.020 ;
  LAYER metal3 ;
  RECT 1444.720 97.780 1445.840 101.020 ;
  LAYER metal2 ;
  RECT 1444.720 97.780 1445.840 101.020 ;
  LAYER metal1 ;
  RECT 1444.720 97.780 1445.840 101.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 89.940 1445.840 93.180 ;
  LAYER metal4 ;
  RECT 1444.720 89.940 1445.840 93.180 ;
  LAYER metal3 ;
  RECT 1444.720 89.940 1445.840 93.180 ;
  LAYER metal2 ;
  RECT 1444.720 89.940 1445.840 93.180 ;
  LAYER metal1 ;
  RECT 1444.720 89.940 1445.840 93.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 50.740 1445.840 53.980 ;
  LAYER metal4 ;
  RECT 1444.720 50.740 1445.840 53.980 ;
  LAYER metal3 ;
  RECT 1444.720 50.740 1445.840 53.980 ;
  LAYER metal2 ;
  RECT 1444.720 50.740 1445.840 53.980 ;
  LAYER metal1 ;
  RECT 1444.720 50.740 1445.840 53.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 42.900 1445.840 46.140 ;
  LAYER metal4 ;
  RECT 1444.720 42.900 1445.840 46.140 ;
  LAYER metal3 ;
  RECT 1444.720 42.900 1445.840 46.140 ;
  LAYER metal2 ;
  RECT 1444.720 42.900 1445.840 46.140 ;
  LAYER metal1 ;
  RECT 1444.720 42.900 1445.840 46.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 35.060 1445.840 38.300 ;
  LAYER metal4 ;
  RECT 1444.720 35.060 1445.840 38.300 ;
  LAYER metal3 ;
  RECT 1444.720 35.060 1445.840 38.300 ;
  LAYER metal2 ;
  RECT 1444.720 35.060 1445.840 38.300 ;
  LAYER metal1 ;
  RECT 1444.720 35.060 1445.840 38.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 27.220 1445.840 30.460 ;
  LAYER metal4 ;
  RECT 1444.720 27.220 1445.840 30.460 ;
  LAYER metal3 ;
  RECT 1444.720 27.220 1445.840 30.460 ;
  LAYER metal2 ;
  RECT 1444.720 27.220 1445.840 30.460 ;
  LAYER metal1 ;
  RECT 1444.720 27.220 1445.840 30.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 19.380 1445.840 22.620 ;
  LAYER metal4 ;
  RECT 1444.720 19.380 1445.840 22.620 ;
  LAYER metal3 ;
  RECT 1444.720 19.380 1445.840 22.620 ;
  LAYER metal2 ;
  RECT 1444.720 19.380 1445.840 22.620 ;
  LAYER metal1 ;
  RECT 1444.720 19.380 1445.840 22.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 11.540 1445.840 14.780 ;
  LAYER metal4 ;
  RECT 1444.720 11.540 1445.840 14.780 ;
  LAYER metal3 ;
  RECT 1444.720 11.540 1445.840 14.780 ;
  LAYER metal2 ;
  RECT 1444.720 11.540 1445.840 14.780 ;
  LAYER metal1 ;
  RECT 1444.720 11.540 1445.840 14.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 521.140 1.120 524.380 ;
  LAYER metal4 ;
  RECT 0.000 521.140 1.120 524.380 ;
  LAYER metal3 ;
  RECT 0.000 521.140 1.120 524.380 ;
  LAYER metal2 ;
  RECT 0.000 521.140 1.120 524.380 ;
  LAYER metal1 ;
  RECT 0.000 521.140 1.120 524.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 513.300 1.120 516.540 ;
  LAYER metal4 ;
  RECT 0.000 513.300 1.120 516.540 ;
  LAYER metal3 ;
  RECT 0.000 513.300 1.120 516.540 ;
  LAYER metal2 ;
  RECT 0.000 513.300 1.120 516.540 ;
  LAYER metal1 ;
  RECT 0.000 513.300 1.120 516.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 505.460 1.120 508.700 ;
  LAYER metal4 ;
  RECT 0.000 505.460 1.120 508.700 ;
  LAYER metal3 ;
  RECT 0.000 505.460 1.120 508.700 ;
  LAYER metal2 ;
  RECT 0.000 505.460 1.120 508.700 ;
  LAYER metal1 ;
  RECT 0.000 505.460 1.120 508.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 497.620 1.120 500.860 ;
  LAYER metal4 ;
  RECT 0.000 497.620 1.120 500.860 ;
  LAYER metal3 ;
  RECT 0.000 497.620 1.120 500.860 ;
  LAYER metal2 ;
  RECT 0.000 497.620 1.120 500.860 ;
  LAYER metal1 ;
  RECT 0.000 497.620 1.120 500.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 489.780 1.120 493.020 ;
  LAYER metal4 ;
  RECT 0.000 489.780 1.120 493.020 ;
  LAYER metal3 ;
  RECT 0.000 489.780 1.120 493.020 ;
  LAYER metal2 ;
  RECT 0.000 489.780 1.120 493.020 ;
  LAYER metal1 ;
  RECT 0.000 489.780 1.120 493.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 481.940 1.120 485.180 ;
  LAYER metal4 ;
  RECT 0.000 481.940 1.120 485.180 ;
  LAYER metal3 ;
  RECT 0.000 481.940 1.120 485.180 ;
  LAYER metal2 ;
  RECT 0.000 481.940 1.120 485.180 ;
  LAYER metal1 ;
  RECT 0.000 481.940 1.120 485.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 442.740 1.120 445.980 ;
  LAYER metal4 ;
  RECT 0.000 442.740 1.120 445.980 ;
  LAYER metal3 ;
  RECT 0.000 442.740 1.120 445.980 ;
  LAYER metal2 ;
  RECT 0.000 442.740 1.120 445.980 ;
  LAYER metal1 ;
  RECT 0.000 442.740 1.120 445.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 434.900 1.120 438.140 ;
  LAYER metal4 ;
  RECT 0.000 434.900 1.120 438.140 ;
  LAYER metal3 ;
  RECT 0.000 434.900 1.120 438.140 ;
  LAYER metal2 ;
  RECT 0.000 434.900 1.120 438.140 ;
  LAYER metal1 ;
  RECT 0.000 434.900 1.120 438.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 427.060 1.120 430.300 ;
  LAYER metal4 ;
  RECT 0.000 427.060 1.120 430.300 ;
  LAYER metal3 ;
  RECT 0.000 427.060 1.120 430.300 ;
  LAYER metal2 ;
  RECT 0.000 427.060 1.120 430.300 ;
  LAYER metal1 ;
  RECT 0.000 427.060 1.120 430.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 419.220 1.120 422.460 ;
  LAYER metal4 ;
  RECT 0.000 419.220 1.120 422.460 ;
  LAYER metal3 ;
  RECT 0.000 419.220 1.120 422.460 ;
  LAYER metal2 ;
  RECT 0.000 419.220 1.120 422.460 ;
  LAYER metal1 ;
  RECT 0.000 419.220 1.120 422.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 411.380 1.120 414.620 ;
  LAYER metal4 ;
  RECT 0.000 411.380 1.120 414.620 ;
  LAYER metal3 ;
  RECT 0.000 411.380 1.120 414.620 ;
  LAYER metal2 ;
  RECT 0.000 411.380 1.120 414.620 ;
  LAYER metal1 ;
  RECT 0.000 411.380 1.120 414.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 403.540 1.120 406.780 ;
  LAYER metal4 ;
  RECT 0.000 403.540 1.120 406.780 ;
  LAYER metal3 ;
  RECT 0.000 403.540 1.120 406.780 ;
  LAYER metal2 ;
  RECT 0.000 403.540 1.120 406.780 ;
  LAYER metal1 ;
  RECT 0.000 403.540 1.120 406.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 364.340 1.120 367.580 ;
  LAYER metal4 ;
  RECT 0.000 364.340 1.120 367.580 ;
  LAYER metal3 ;
  RECT 0.000 364.340 1.120 367.580 ;
  LAYER metal2 ;
  RECT 0.000 364.340 1.120 367.580 ;
  LAYER metal1 ;
  RECT 0.000 364.340 1.120 367.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 356.500 1.120 359.740 ;
  LAYER metal4 ;
  RECT 0.000 356.500 1.120 359.740 ;
  LAYER metal3 ;
  RECT 0.000 356.500 1.120 359.740 ;
  LAYER metal2 ;
  RECT 0.000 356.500 1.120 359.740 ;
  LAYER metal1 ;
  RECT 0.000 356.500 1.120 359.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 348.660 1.120 351.900 ;
  LAYER metal4 ;
  RECT 0.000 348.660 1.120 351.900 ;
  LAYER metal3 ;
  RECT 0.000 348.660 1.120 351.900 ;
  LAYER metal2 ;
  RECT 0.000 348.660 1.120 351.900 ;
  LAYER metal1 ;
  RECT 0.000 348.660 1.120 351.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 340.820 1.120 344.060 ;
  LAYER metal4 ;
  RECT 0.000 340.820 1.120 344.060 ;
  LAYER metal3 ;
  RECT 0.000 340.820 1.120 344.060 ;
  LAYER metal2 ;
  RECT 0.000 340.820 1.120 344.060 ;
  LAYER metal1 ;
  RECT 0.000 340.820 1.120 344.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 332.980 1.120 336.220 ;
  LAYER metal4 ;
  RECT 0.000 332.980 1.120 336.220 ;
  LAYER metal3 ;
  RECT 0.000 332.980 1.120 336.220 ;
  LAYER metal2 ;
  RECT 0.000 332.980 1.120 336.220 ;
  LAYER metal1 ;
  RECT 0.000 332.980 1.120 336.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 325.140 1.120 328.380 ;
  LAYER metal4 ;
  RECT 0.000 325.140 1.120 328.380 ;
  LAYER metal3 ;
  RECT 0.000 325.140 1.120 328.380 ;
  LAYER metal2 ;
  RECT 0.000 325.140 1.120 328.380 ;
  LAYER metal1 ;
  RECT 0.000 325.140 1.120 328.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 285.940 1.120 289.180 ;
  LAYER metal4 ;
  RECT 0.000 285.940 1.120 289.180 ;
  LAYER metal3 ;
  RECT 0.000 285.940 1.120 289.180 ;
  LAYER metal2 ;
  RECT 0.000 285.940 1.120 289.180 ;
  LAYER metal1 ;
  RECT 0.000 285.940 1.120 289.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 278.100 1.120 281.340 ;
  LAYER metal4 ;
  RECT 0.000 278.100 1.120 281.340 ;
  LAYER metal3 ;
  RECT 0.000 278.100 1.120 281.340 ;
  LAYER metal2 ;
  RECT 0.000 278.100 1.120 281.340 ;
  LAYER metal1 ;
  RECT 0.000 278.100 1.120 281.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 270.260 1.120 273.500 ;
  LAYER metal4 ;
  RECT 0.000 270.260 1.120 273.500 ;
  LAYER metal3 ;
  RECT 0.000 270.260 1.120 273.500 ;
  LAYER metal2 ;
  RECT 0.000 270.260 1.120 273.500 ;
  LAYER metal1 ;
  RECT 0.000 270.260 1.120 273.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 262.420 1.120 265.660 ;
  LAYER metal4 ;
  RECT 0.000 262.420 1.120 265.660 ;
  LAYER metal3 ;
  RECT 0.000 262.420 1.120 265.660 ;
  LAYER metal2 ;
  RECT 0.000 262.420 1.120 265.660 ;
  LAYER metal1 ;
  RECT 0.000 262.420 1.120 265.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 254.580 1.120 257.820 ;
  LAYER metal4 ;
  RECT 0.000 254.580 1.120 257.820 ;
  LAYER metal3 ;
  RECT 0.000 254.580 1.120 257.820 ;
  LAYER metal2 ;
  RECT 0.000 254.580 1.120 257.820 ;
  LAYER metal1 ;
  RECT 0.000 254.580 1.120 257.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 246.740 1.120 249.980 ;
  LAYER metal4 ;
  RECT 0.000 246.740 1.120 249.980 ;
  LAYER metal3 ;
  RECT 0.000 246.740 1.120 249.980 ;
  LAYER metal2 ;
  RECT 0.000 246.740 1.120 249.980 ;
  LAYER metal1 ;
  RECT 0.000 246.740 1.120 249.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 207.540 1.120 210.780 ;
  LAYER metal4 ;
  RECT 0.000 207.540 1.120 210.780 ;
  LAYER metal3 ;
  RECT 0.000 207.540 1.120 210.780 ;
  LAYER metal2 ;
  RECT 0.000 207.540 1.120 210.780 ;
  LAYER metal1 ;
  RECT 0.000 207.540 1.120 210.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER metal4 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER metal3 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER metal2 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER metal1 ;
  RECT 0.000 199.700 1.120 202.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER metal4 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER metal3 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER metal2 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER metal1 ;
  RECT 0.000 191.860 1.120 195.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER metal4 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER metal3 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER metal2 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER metal1 ;
  RECT 0.000 184.020 1.120 187.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER metal4 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER metal3 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER metal2 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER metal1 ;
  RECT 0.000 176.180 1.120 179.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER metal4 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER metal3 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER metal2 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER metal1 ;
  RECT 0.000 168.340 1.120 171.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER metal4 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER metal3 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER metal2 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER metal1 ;
  RECT 0.000 129.140 1.120 132.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER metal4 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER metal3 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER metal2 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER metal1 ;
  RECT 0.000 121.300 1.120 124.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER metal4 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER metal3 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER metal2 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER metal1 ;
  RECT 0.000 113.460 1.120 116.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER metal4 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER metal3 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER metal2 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER metal1 ;
  RECT 0.000 105.620 1.120 108.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER metal4 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER metal3 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER metal2 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER metal1 ;
  RECT 0.000 97.780 1.120 101.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER metal4 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER metal3 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER metal2 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER metal1 ;
  RECT 0.000 89.940 1.120 93.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER metal4 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER metal3 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER metal2 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER metal1 ;
  RECT 0.000 50.740 1.120 53.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER metal4 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER metal3 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER metal2 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER metal1 ;
  RECT 0.000 42.900 1.120 46.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER metal4 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER metal3 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER metal2 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER metal1 ;
  RECT 0.000 35.060 1.120 38.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER metal4 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER metal3 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER metal2 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER metal1 ;
  RECT 0.000 27.220 1.120 30.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER metal4 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER metal3 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER metal2 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER metal1 ;
  RECT 0.000 19.380 1.120 22.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER metal4 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER metal3 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER metal2 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER metal1 ;
  RECT 0.000 11.540 1.120 14.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1433.840 543.200 1437.380 544.320 ;
  LAYER metal4 ;
  RECT 1433.840 543.200 1437.380 544.320 ;
  LAYER metal3 ;
  RECT 1433.840 543.200 1437.380 544.320 ;
  LAYER metal2 ;
  RECT 1433.840 543.200 1437.380 544.320 ;
  LAYER metal1 ;
  RECT 1433.840 543.200 1437.380 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1425.160 543.200 1428.700 544.320 ;
  LAYER metal4 ;
  RECT 1425.160 543.200 1428.700 544.320 ;
  LAYER metal3 ;
  RECT 1425.160 543.200 1428.700 544.320 ;
  LAYER metal2 ;
  RECT 1425.160 543.200 1428.700 544.320 ;
  LAYER metal1 ;
  RECT 1425.160 543.200 1428.700 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1411.520 543.200 1415.060 544.320 ;
  LAYER metal4 ;
  RECT 1411.520 543.200 1415.060 544.320 ;
  LAYER metal3 ;
  RECT 1411.520 543.200 1415.060 544.320 ;
  LAYER metal2 ;
  RECT 1411.520 543.200 1415.060 544.320 ;
  LAYER metal1 ;
  RECT 1411.520 543.200 1415.060 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1397.880 543.200 1401.420 544.320 ;
  LAYER metal4 ;
  RECT 1397.880 543.200 1401.420 544.320 ;
  LAYER metal3 ;
  RECT 1397.880 543.200 1401.420 544.320 ;
  LAYER metal2 ;
  RECT 1397.880 543.200 1401.420 544.320 ;
  LAYER metal1 ;
  RECT 1397.880 543.200 1401.420 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1384.860 543.200 1388.400 544.320 ;
  LAYER metal4 ;
  RECT 1384.860 543.200 1388.400 544.320 ;
  LAYER metal3 ;
  RECT 1384.860 543.200 1388.400 544.320 ;
  LAYER metal2 ;
  RECT 1384.860 543.200 1388.400 544.320 ;
  LAYER metal1 ;
  RECT 1384.860 543.200 1388.400 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1371.220 543.200 1374.760 544.320 ;
  LAYER metal4 ;
  RECT 1371.220 543.200 1374.760 544.320 ;
  LAYER metal3 ;
  RECT 1371.220 543.200 1374.760 544.320 ;
  LAYER metal2 ;
  RECT 1371.220 543.200 1374.760 544.320 ;
  LAYER metal1 ;
  RECT 1371.220 543.200 1374.760 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1304.260 543.200 1307.800 544.320 ;
  LAYER metal4 ;
  RECT 1304.260 543.200 1307.800 544.320 ;
  LAYER metal3 ;
  RECT 1304.260 543.200 1307.800 544.320 ;
  LAYER metal2 ;
  RECT 1304.260 543.200 1307.800 544.320 ;
  LAYER metal1 ;
  RECT 1304.260 543.200 1307.800 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1290.620 543.200 1294.160 544.320 ;
  LAYER metal4 ;
  RECT 1290.620 543.200 1294.160 544.320 ;
  LAYER metal3 ;
  RECT 1290.620 543.200 1294.160 544.320 ;
  LAYER metal2 ;
  RECT 1290.620 543.200 1294.160 544.320 ;
  LAYER metal1 ;
  RECT 1290.620 543.200 1294.160 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1276.980 543.200 1280.520 544.320 ;
  LAYER metal4 ;
  RECT 1276.980 543.200 1280.520 544.320 ;
  LAYER metal3 ;
  RECT 1276.980 543.200 1280.520 544.320 ;
  LAYER metal2 ;
  RECT 1276.980 543.200 1280.520 544.320 ;
  LAYER metal1 ;
  RECT 1276.980 543.200 1280.520 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1263.960 543.200 1267.500 544.320 ;
  LAYER metal4 ;
  RECT 1263.960 543.200 1267.500 544.320 ;
  LAYER metal3 ;
  RECT 1263.960 543.200 1267.500 544.320 ;
  LAYER metal2 ;
  RECT 1263.960 543.200 1267.500 544.320 ;
  LAYER metal1 ;
  RECT 1263.960 543.200 1267.500 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1250.320 543.200 1253.860 544.320 ;
  LAYER metal4 ;
  RECT 1250.320 543.200 1253.860 544.320 ;
  LAYER metal3 ;
  RECT 1250.320 543.200 1253.860 544.320 ;
  LAYER metal2 ;
  RECT 1250.320 543.200 1253.860 544.320 ;
  LAYER metal1 ;
  RECT 1250.320 543.200 1253.860 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1236.680 543.200 1240.220 544.320 ;
  LAYER metal4 ;
  RECT 1236.680 543.200 1240.220 544.320 ;
  LAYER metal3 ;
  RECT 1236.680 543.200 1240.220 544.320 ;
  LAYER metal2 ;
  RECT 1236.680 543.200 1240.220 544.320 ;
  LAYER metal1 ;
  RECT 1236.680 543.200 1240.220 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1169.720 543.200 1173.260 544.320 ;
  LAYER metal4 ;
  RECT 1169.720 543.200 1173.260 544.320 ;
  LAYER metal3 ;
  RECT 1169.720 543.200 1173.260 544.320 ;
  LAYER metal2 ;
  RECT 1169.720 543.200 1173.260 544.320 ;
  LAYER metal1 ;
  RECT 1169.720 543.200 1173.260 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1156.080 543.200 1159.620 544.320 ;
  LAYER metal4 ;
  RECT 1156.080 543.200 1159.620 544.320 ;
  LAYER metal3 ;
  RECT 1156.080 543.200 1159.620 544.320 ;
  LAYER metal2 ;
  RECT 1156.080 543.200 1159.620 544.320 ;
  LAYER metal1 ;
  RECT 1156.080 543.200 1159.620 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1143.060 543.200 1146.600 544.320 ;
  LAYER metal4 ;
  RECT 1143.060 543.200 1146.600 544.320 ;
  LAYER metal3 ;
  RECT 1143.060 543.200 1146.600 544.320 ;
  LAYER metal2 ;
  RECT 1143.060 543.200 1146.600 544.320 ;
  LAYER metal1 ;
  RECT 1143.060 543.200 1146.600 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1129.420 543.200 1132.960 544.320 ;
  LAYER metal4 ;
  RECT 1129.420 543.200 1132.960 544.320 ;
  LAYER metal3 ;
  RECT 1129.420 543.200 1132.960 544.320 ;
  LAYER metal2 ;
  RECT 1129.420 543.200 1132.960 544.320 ;
  LAYER metal1 ;
  RECT 1129.420 543.200 1132.960 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1115.780 543.200 1119.320 544.320 ;
  LAYER metal4 ;
  RECT 1115.780 543.200 1119.320 544.320 ;
  LAYER metal3 ;
  RECT 1115.780 543.200 1119.320 544.320 ;
  LAYER metal2 ;
  RECT 1115.780 543.200 1119.320 544.320 ;
  LAYER metal1 ;
  RECT 1115.780 543.200 1119.320 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1102.760 543.200 1106.300 544.320 ;
  LAYER metal4 ;
  RECT 1102.760 543.200 1106.300 544.320 ;
  LAYER metal3 ;
  RECT 1102.760 543.200 1106.300 544.320 ;
  LAYER metal2 ;
  RECT 1102.760 543.200 1106.300 544.320 ;
  LAYER metal1 ;
  RECT 1102.760 543.200 1106.300 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1035.180 543.200 1038.720 544.320 ;
  LAYER metal4 ;
  RECT 1035.180 543.200 1038.720 544.320 ;
  LAYER metal3 ;
  RECT 1035.180 543.200 1038.720 544.320 ;
  LAYER metal2 ;
  RECT 1035.180 543.200 1038.720 544.320 ;
  LAYER metal1 ;
  RECT 1035.180 543.200 1038.720 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1021.540 543.200 1025.080 544.320 ;
  LAYER metal4 ;
  RECT 1021.540 543.200 1025.080 544.320 ;
  LAYER metal3 ;
  RECT 1021.540 543.200 1025.080 544.320 ;
  LAYER metal2 ;
  RECT 1021.540 543.200 1025.080 544.320 ;
  LAYER metal1 ;
  RECT 1021.540 543.200 1025.080 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1010.380 543.200 1013.920 544.320 ;
  LAYER metal4 ;
  RECT 1010.380 543.200 1013.920 544.320 ;
  LAYER metal3 ;
  RECT 1010.380 543.200 1013.920 544.320 ;
  LAYER metal2 ;
  RECT 1010.380 543.200 1013.920 544.320 ;
  LAYER metal1 ;
  RECT 1010.380 543.200 1013.920 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 994.880 543.200 998.420 544.320 ;
  LAYER metal4 ;
  RECT 994.880 543.200 998.420 544.320 ;
  LAYER metal3 ;
  RECT 994.880 543.200 998.420 544.320 ;
  LAYER metal2 ;
  RECT 994.880 543.200 998.420 544.320 ;
  LAYER metal1 ;
  RECT 994.880 543.200 998.420 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 981.240 543.200 984.780 544.320 ;
  LAYER metal4 ;
  RECT 981.240 543.200 984.780 544.320 ;
  LAYER metal3 ;
  RECT 981.240 543.200 984.780 544.320 ;
  LAYER metal2 ;
  RECT 981.240 543.200 984.780 544.320 ;
  LAYER metal1 ;
  RECT 981.240 543.200 984.780 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 968.220 543.200 971.760 544.320 ;
  LAYER metal4 ;
  RECT 968.220 543.200 971.760 544.320 ;
  LAYER metal3 ;
  RECT 968.220 543.200 971.760 544.320 ;
  LAYER metal2 ;
  RECT 968.220 543.200 971.760 544.320 ;
  LAYER metal1 ;
  RECT 968.220 543.200 971.760 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 900.640 543.200 904.180 544.320 ;
  LAYER metal4 ;
  RECT 900.640 543.200 904.180 544.320 ;
  LAYER metal3 ;
  RECT 900.640 543.200 904.180 544.320 ;
  LAYER metal2 ;
  RECT 900.640 543.200 904.180 544.320 ;
  LAYER metal1 ;
  RECT 900.640 543.200 904.180 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 887.620 543.200 891.160 544.320 ;
  LAYER metal4 ;
  RECT 887.620 543.200 891.160 544.320 ;
  LAYER metal3 ;
  RECT 887.620 543.200 891.160 544.320 ;
  LAYER metal2 ;
  RECT 887.620 543.200 891.160 544.320 ;
  LAYER metal1 ;
  RECT 887.620 543.200 891.160 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 873.980 543.200 877.520 544.320 ;
  LAYER metal4 ;
  RECT 873.980 543.200 877.520 544.320 ;
  LAYER metal3 ;
  RECT 873.980 543.200 877.520 544.320 ;
  LAYER metal2 ;
  RECT 873.980 543.200 877.520 544.320 ;
  LAYER metal1 ;
  RECT 873.980 543.200 877.520 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 860.340 543.200 863.880 544.320 ;
  LAYER metal4 ;
  RECT 860.340 543.200 863.880 544.320 ;
  LAYER metal3 ;
  RECT 860.340 543.200 863.880 544.320 ;
  LAYER metal2 ;
  RECT 860.340 543.200 863.880 544.320 ;
  LAYER metal1 ;
  RECT 860.340 543.200 863.880 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 847.320 543.200 850.860 544.320 ;
  LAYER metal4 ;
  RECT 847.320 543.200 850.860 544.320 ;
  LAYER metal3 ;
  RECT 847.320 543.200 850.860 544.320 ;
  LAYER metal2 ;
  RECT 847.320 543.200 850.860 544.320 ;
  LAYER metal1 ;
  RECT 847.320 543.200 850.860 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 833.680 543.200 837.220 544.320 ;
  LAYER metal4 ;
  RECT 833.680 543.200 837.220 544.320 ;
  LAYER metal3 ;
  RECT 833.680 543.200 837.220 544.320 ;
  LAYER metal2 ;
  RECT 833.680 543.200 837.220 544.320 ;
  LAYER metal1 ;
  RECT 833.680 543.200 837.220 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 766.720 543.200 770.260 544.320 ;
  LAYER metal4 ;
  RECT 766.720 543.200 770.260 544.320 ;
  LAYER metal3 ;
  RECT 766.720 543.200 770.260 544.320 ;
  LAYER metal2 ;
  RECT 766.720 543.200 770.260 544.320 ;
  LAYER metal1 ;
  RECT 766.720 543.200 770.260 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 753.080 543.200 756.620 544.320 ;
  LAYER metal4 ;
  RECT 753.080 543.200 756.620 544.320 ;
  LAYER metal3 ;
  RECT 753.080 543.200 756.620 544.320 ;
  LAYER metal2 ;
  RECT 753.080 543.200 756.620 544.320 ;
  LAYER metal1 ;
  RECT 753.080 543.200 756.620 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 739.440 543.200 742.980 544.320 ;
  LAYER metal4 ;
  RECT 739.440 543.200 742.980 544.320 ;
  LAYER metal3 ;
  RECT 739.440 543.200 742.980 544.320 ;
  LAYER metal2 ;
  RECT 739.440 543.200 742.980 544.320 ;
  LAYER metal1 ;
  RECT 739.440 543.200 742.980 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 726.420 543.200 729.960 544.320 ;
  LAYER metal4 ;
  RECT 726.420 543.200 729.960 544.320 ;
  LAYER metal3 ;
  RECT 726.420 543.200 729.960 544.320 ;
  LAYER metal2 ;
  RECT 726.420 543.200 729.960 544.320 ;
  LAYER metal1 ;
  RECT 726.420 543.200 729.960 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 712.780 543.200 716.320 544.320 ;
  LAYER metal4 ;
  RECT 712.780 543.200 716.320 544.320 ;
  LAYER metal3 ;
  RECT 712.780 543.200 716.320 544.320 ;
  LAYER metal2 ;
  RECT 712.780 543.200 716.320 544.320 ;
  LAYER metal1 ;
  RECT 712.780 543.200 716.320 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 699.140 543.200 702.680 544.320 ;
  LAYER metal4 ;
  RECT 699.140 543.200 702.680 544.320 ;
  LAYER metal3 ;
  RECT 699.140 543.200 702.680 544.320 ;
  LAYER metal2 ;
  RECT 699.140 543.200 702.680 544.320 ;
  LAYER metal1 ;
  RECT 699.140 543.200 702.680 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 632.180 543.200 635.720 544.320 ;
  LAYER metal4 ;
  RECT 632.180 543.200 635.720 544.320 ;
  LAYER metal3 ;
  RECT 632.180 543.200 635.720 544.320 ;
  LAYER metal2 ;
  RECT 632.180 543.200 635.720 544.320 ;
  LAYER metal1 ;
  RECT 632.180 543.200 635.720 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 618.540 543.200 622.080 544.320 ;
  LAYER metal4 ;
  RECT 618.540 543.200 622.080 544.320 ;
  LAYER metal3 ;
  RECT 618.540 543.200 622.080 544.320 ;
  LAYER metal2 ;
  RECT 618.540 543.200 622.080 544.320 ;
  LAYER metal1 ;
  RECT 618.540 543.200 622.080 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 604.900 543.200 608.440 544.320 ;
  LAYER metal4 ;
  RECT 604.900 543.200 608.440 544.320 ;
  LAYER metal3 ;
  RECT 604.900 543.200 608.440 544.320 ;
  LAYER metal2 ;
  RECT 604.900 543.200 608.440 544.320 ;
  LAYER metal1 ;
  RECT 604.900 543.200 608.440 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 591.880 543.200 595.420 544.320 ;
  LAYER metal4 ;
  RECT 591.880 543.200 595.420 544.320 ;
  LAYER metal3 ;
  RECT 591.880 543.200 595.420 544.320 ;
  LAYER metal2 ;
  RECT 591.880 543.200 595.420 544.320 ;
  LAYER metal1 ;
  RECT 591.880 543.200 595.420 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 580.720 543.200 584.260 544.320 ;
  LAYER metal4 ;
  RECT 580.720 543.200 584.260 544.320 ;
  LAYER metal3 ;
  RECT 580.720 543.200 584.260 544.320 ;
  LAYER metal2 ;
  RECT 580.720 543.200 584.260 544.320 ;
  LAYER metal1 ;
  RECT 580.720 543.200 584.260 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 564.600 543.200 568.140 544.320 ;
  LAYER metal4 ;
  RECT 564.600 543.200 568.140 544.320 ;
  LAYER metal3 ;
  RECT 564.600 543.200 568.140 544.320 ;
  LAYER metal2 ;
  RECT 564.600 543.200 568.140 544.320 ;
  LAYER metal1 ;
  RECT 564.600 543.200 568.140 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 470.980 543.200 474.520 544.320 ;
  LAYER metal4 ;
  RECT 470.980 543.200 474.520 544.320 ;
  LAYER metal3 ;
  RECT 470.980 543.200 474.520 544.320 ;
  LAYER metal2 ;
  RECT 470.980 543.200 474.520 544.320 ;
  LAYER metal1 ;
  RECT 470.980 543.200 474.520 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 462.300 543.200 465.840 544.320 ;
  LAYER metal4 ;
  RECT 462.300 543.200 465.840 544.320 ;
  LAYER metal3 ;
  RECT 462.300 543.200 465.840 544.320 ;
  LAYER metal2 ;
  RECT 462.300 543.200 465.840 544.320 ;
  LAYER metal1 ;
  RECT 462.300 543.200 465.840 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 453.620 543.200 457.160 544.320 ;
  LAYER metal4 ;
  RECT 453.620 543.200 457.160 544.320 ;
  LAYER metal3 ;
  RECT 453.620 543.200 457.160 544.320 ;
  LAYER metal2 ;
  RECT 453.620 543.200 457.160 544.320 ;
  LAYER metal1 ;
  RECT 453.620 543.200 457.160 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 439.980 543.200 443.520 544.320 ;
  LAYER metal4 ;
  RECT 439.980 543.200 443.520 544.320 ;
  LAYER metal3 ;
  RECT 439.980 543.200 443.520 544.320 ;
  LAYER metal2 ;
  RECT 439.980 543.200 443.520 544.320 ;
  LAYER metal1 ;
  RECT 439.980 543.200 443.520 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 431.300 543.200 434.840 544.320 ;
  LAYER metal4 ;
  RECT 431.300 543.200 434.840 544.320 ;
  LAYER metal3 ;
  RECT 431.300 543.200 434.840 544.320 ;
  LAYER metal2 ;
  RECT 431.300 543.200 434.840 544.320 ;
  LAYER metal1 ;
  RECT 431.300 543.200 434.840 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 418.280 543.200 421.820 544.320 ;
  LAYER metal4 ;
  RECT 418.280 543.200 421.820 544.320 ;
  LAYER metal3 ;
  RECT 418.280 543.200 421.820 544.320 ;
  LAYER metal2 ;
  RECT 418.280 543.200 421.820 544.320 ;
  LAYER metal1 ;
  RECT 418.280 543.200 421.820 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 350.700 543.200 354.240 544.320 ;
  LAYER metal4 ;
  RECT 350.700 543.200 354.240 544.320 ;
  LAYER metal3 ;
  RECT 350.700 543.200 354.240 544.320 ;
  LAYER metal2 ;
  RECT 350.700 543.200 354.240 544.320 ;
  LAYER metal1 ;
  RECT 350.700 543.200 354.240 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 337.680 543.200 341.220 544.320 ;
  LAYER metal4 ;
  RECT 337.680 543.200 341.220 544.320 ;
  LAYER metal3 ;
  RECT 337.680 543.200 341.220 544.320 ;
  LAYER metal2 ;
  RECT 337.680 543.200 341.220 544.320 ;
  LAYER metal1 ;
  RECT 337.680 543.200 341.220 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 324.040 543.200 327.580 544.320 ;
  LAYER metal4 ;
  RECT 324.040 543.200 327.580 544.320 ;
  LAYER metal3 ;
  RECT 324.040 543.200 327.580 544.320 ;
  LAYER metal2 ;
  RECT 324.040 543.200 327.580 544.320 ;
  LAYER metal1 ;
  RECT 324.040 543.200 327.580 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 310.400 543.200 313.940 544.320 ;
  LAYER metal4 ;
  RECT 310.400 543.200 313.940 544.320 ;
  LAYER metal3 ;
  RECT 310.400 543.200 313.940 544.320 ;
  LAYER metal2 ;
  RECT 310.400 543.200 313.940 544.320 ;
  LAYER metal1 ;
  RECT 310.400 543.200 313.940 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 297.380 543.200 300.920 544.320 ;
  LAYER metal4 ;
  RECT 297.380 543.200 300.920 544.320 ;
  LAYER metal3 ;
  RECT 297.380 543.200 300.920 544.320 ;
  LAYER metal2 ;
  RECT 297.380 543.200 300.920 544.320 ;
  LAYER metal1 ;
  RECT 297.380 543.200 300.920 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 283.740 543.200 287.280 544.320 ;
  LAYER metal4 ;
  RECT 283.740 543.200 287.280 544.320 ;
  LAYER metal3 ;
  RECT 283.740 543.200 287.280 544.320 ;
  LAYER metal2 ;
  RECT 283.740 543.200 287.280 544.320 ;
  LAYER metal1 ;
  RECT 283.740 543.200 287.280 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 216.780 543.200 220.320 544.320 ;
  LAYER metal4 ;
  RECT 216.780 543.200 220.320 544.320 ;
  LAYER metal3 ;
  RECT 216.780 543.200 220.320 544.320 ;
  LAYER metal2 ;
  RECT 216.780 543.200 220.320 544.320 ;
  LAYER metal1 ;
  RECT 216.780 543.200 220.320 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 203.140 543.200 206.680 544.320 ;
  LAYER metal4 ;
  RECT 203.140 543.200 206.680 544.320 ;
  LAYER metal3 ;
  RECT 203.140 543.200 206.680 544.320 ;
  LAYER metal2 ;
  RECT 203.140 543.200 206.680 544.320 ;
  LAYER metal1 ;
  RECT 203.140 543.200 206.680 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 189.500 543.200 193.040 544.320 ;
  LAYER metal4 ;
  RECT 189.500 543.200 193.040 544.320 ;
  LAYER metal3 ;
  RECT 189.500 543.200 193.040 544.320 ;
  LAYER metal2 ;
  RECT 189.500 543.200 193.040 544.320 ;
  LAYER metal1 ;
  RECT 189.500 543.200 193.040 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 176.480 543.200 180.020 544.320 ;
  LAYER metal4 ;
  RECT 176.480 543.200 180.020 544.320 ;
  LAYER metal3 ;
  RECT 176.480 543.200 180.020 544.320 ;
  LAYER metal2 ;
  RECT 176.480 543.200 180.020 544.320 ;
  LAYER metal1 ;
  RECT 176.480 543.200 180.020 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 162.840 543.200 166.380 544.320 ;
  LAYER metal4 ;
  RECT 162.840 543.200 166.380 544.320 ;
  LAYER metal3 ;
  RECT 162.840 543.200 166.380 544.320 ;
  LAYER metal2 ;
  RECT 162.840 543.200 166.380 544.320 ;
  LAYER metal1 ;
  RECT 162.840 543.200 166.380 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 149.200 543.200 152.740 544.320 ;
  LAYER metal4 ;
  RECT 149.200 543.200 152.740 544.320 ;
  LAYER metal3 ;
  RECT 149.200 543.200 152.740 544.320 ;
  LAYER metal2 ;
  RECT 149.200 543.200 152.740 544.320 ;
  LAYER metal1 ;
  RECT 149.200 543.200 152.740 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 82.240 543.200 85.780 544.320 ;
  LAYER metal4 ;
  RECT 82.240 543.200 85.780 544.320 ;
  LAYER metal3 ;
  RECT 82.240 543.200 85.780 544.320 ;
  LAYER metal2 ;
  RECT 82.240 543.200 85.780 544.320 ;
  LAYER metal1 ;
  RECT 82.240 543.200 85.780 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 68.600 543.200 72.140 544.320 ;
  LAYER metal4 ;
  RECT 68.600 543.200 72.140 544.320 ;
  LAYER metal3 ;
  RECT 68.600 543.200 72.140 544.320 ;
  LAYER metal2 ;
  RECT 68.600 543.200 72.140 544.320 ;
  LAYER metal1 ;
  RECT 68.600 543.200 72.140 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 54.960 543.200 58.500 544.320 ;
  LAYER metal4 ;
  RECT 54.960 543.200 58.500 544.320 ;
  LAYER metal3 ;
  RECT 54.960 543.200 58.500 544.320 ;
  LAYER metal2 ;
  RECT 54.960 543.200 58.500 544.320 ;
  LAYER metal1 ;
  RECT 54.960 543.200 58.500 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 41.940 543.200 45.480 544.320 ;
  LAYER metal4 ;
  RECT 41.940 543.200 45.480 544.320 ;
  LAYER metal3 ;
  RECT 41.940 543.200 45.480 544.320 ;
  LAYER metal2 ;
  RECT 41.940 543.200 45.480 544.320 ;
  LAYER metal1 ;
  RECT 41.940 543.200 45.480 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 28.300 543.200 31.840 544.320 ;
  LAYER metal4 ;
  RECT 28.300 543.200 31.840 544.320 ;
  LAYER metal3 ;
  RECT 28.300 543.200 31.840 544.320 ;
  LAYER metal2 ;
  RECT 28.300 543.200 31.840 544.320 ;
  LAYER metal1 ;
  RECT 28.300 543.200 31.840 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 17.140 543.200 20.680 544.320 ;
  LAYER metal4 ;
  RECT 17.140 543.200 20.680 544.320 ;
  LAYER metal3 ;
  RECT 17.140 543.200 20.680 544.320 ;
  LAYER metal2 ;
  RECT 17.140 543.200 20.680 544.320 ;
  LAYER metal1 ;
  RECT 17.140 543.200 20.680 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1433.840 0.000 1437.380 1.120 ;
  LAYER metal4 ;
  RECT 1433.840 0.000 1437.380 1.120 ;
  LAYER metal3 ;
  RECT 1433.840 0.000 1437.380 1.120 ;
  LAYER metal2 ;
  RECT 1433.840 0.000 1437.380 1.120 ;
  LAYER metal1 ;
  RECT 1433.840 0.000 1437.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1425.160 0.000 1428.700 1.120 ;
  LAYER metal4 ;
  RECT 1425.160 0.000 1428.700 1.120 ;
  LAYER metal3 ;
  RECT 1425.160 0.000 1428.700 1.120 ;
  LAYER metal2 ;
  RECT 1425.160 0.000 1428.700 1.120 ;
  LAYER metal1 ;
  RECT 1425.160 0.000 1428.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1411.520 0.000 1415.060 1.120 ;
  LAYER metal4 ;
  RECT 1411.520 0.000 1415.060 1.120 ;
  LAYER metal3 ;
  RECT 1411.520 0.000 1415.060 1.120 ;
  LAYER metal2 ;
  RECT 1411.520 0.000 1415.060 1.120 ;
  LAYER metal1 ;
  RECT 1411.520 0.000 1415.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1397.880 0.000 1401.420 1.120 ;
  LAYER metal4 ;
  RECT 1397.880 0.000 1401.420 1.120 ;
  LAYER metal3 ;
  RECT 1397.880 0.000 1401.420 1.120 ;
  LAYER metal2 ;
  RECT 1397.880 0.000 1401.420 1.120 ;
  LAYER metal1 ;
  RECT 1397.880 0.000 1401.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1384.860 0.000 1388.400 1.120 ;
  LAYER metal4 ;
  RECT 1384.860 0.000 1388.400 1.120 ;
  LAYER metal3 ;
  RECT 1384.860 0.000 1388.400 1.120 ;
  LAYER metal2 ;
  RECT 1384.860 0.000 1388.400 1.120 ;
  LAYER metal1 ;
  RECT 1384.860 0.000 1388.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1371.220 0.000 1374.760 1.120 ;
  LAYER metal4 ;
  RECT 1371.220 0.000 1374.760 1.120 ;
  LAYER metal3 ;
  RECT 1371.220 0.000 1374.760 1.120 ;
  LAYER metal2 ;
  RECT 1371.220 0.000 1374.760 1.120 ;
  LAYER metal1 ;
  RECT 1371.220 0.000 1374.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1304.260 0.000 1307.800 1.120 ;
  LAYER metal4 ;
  RECT 1304.260 0.000 1307.800 1.120 ;
  LAYER metal3 ;
  RECT 1304.260 0.000 1307.800 1.120 ;
  LAYER metal2 ;
  RECT 1304.260 0.000 1307.800 1.120 ;
  LAYER metal1 ;
  RECT 1304.260 0.000 1307.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1290.620 0.000 1294.160 1.120 ;
  LAYER metal4 ;
  RECT 1290.620 0.000 1294.160 1.120 ;
  LAYER metal3 ;
  RECT 1290.620 0.000 1294.160 1.120 ;
  LAYER metal2 ;
  RECT 1290.620 0.000 1294.160 1.120 ;
  LAYER metal1 ;
  RECT 1290.620 0.000 1294.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1276.980 0.000 1280.520 1.120 ;
  LAYER metal4 ;
  RECT 1276.980 0.000 1280.520 1.120 ;
  LAYER metal3 ;
  RECT 1276.980 0.000 1280.520 1.120 ;
  LAYER metal2 ;
  RECT 1276.980 0.000 1280.520 1.120 ;
  LAYER metal1 ;
  RECT 1276.980 0.000 1280.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1263.960 0.000 1267.500 1.120 ;
  LAYER metal4 ;
  RECT 1263.960 0.000 1267.500 1.120 ;
  LAYER metal3 ;
  RECT 1263.960 0.000 1267.500 1.120 ;
  LAYER metal2 ;
  RECT 1263.960 0.000 1267.500 1.120 ;
  LAYER metal1 ;
  RECT 1263.960 0.000 1267.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1250.320 0.000 1253.860 1.120 ;
  LAYER metal4 ;
  RECT 1250.320 0.000 1253.860 1.120 ;
  LAYER metal3 ;
  RECT 1250.320 0.000 1253.860 1.120 ;
  LAYER metal2 ;
  RECT 1250.320 0.000 1253.860 1.120 ;
  LAYER metal1 ;
  RECT 1250.320 0.000 1253.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1236.680 0.000 1240.220 1.120 ;
  LAYER metal4 ;
  RECT 1236.680 0.000 1240.220 1.120 ;
  LAYER metal3 ;
  RECT 1236.680 0.000 1240.220 1.120 ;
  LAYER metal2 ;
  RECT 1236.680 0.000 1240.220 1.120 ;
  LAYER metal1 ;
  RECT 1236.680 0.000 1240.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1169.720 0.000 1173.260 1.120 ;
  LAYER metal4 ;
  RECT 1169.720 0.000 1173.260 1.120 ;
  LAYER metal3 ;
  RECT 1169.720 0.000 1173.260 1.120 ;
  LAYER metal2 ;
  RECT 1169.720 0.000 1173.260 1.120 ;
  LAYER metal1 ;
  RECT 1169.720 0.000 1173.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1156.080 0.000 1159.620 1.120 ;
  LAYER metal4 ;
  RECT 1156.080 0.000 1159.620 1.120 ;
  LAYER metal3 ;
  RECT 1156.080 0.000 1159.620 1.120 ;
  LAYER metal2 ;
  RECT 1156.080 0.000 1159.620 1.120 ;
  LAYER metal1 ;
  RECT 1156.080 0.000 1159.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1143.060 0.000 1146.600 1.120 ;
  LAYER metal4 ;
  RECT 1143.060 0.000 1146.600 1.120 ;
  LAYER metal3 ;
  RECT 1143.060 0.000 1146.600 1.120 ;
  LAYER metal2 ;
  RECT 1143.060 0.000 1146.600 1.120 ;
  LAYER metal1 ;
  RECT 1143.060 0.000 1146.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1129.420 0.000 1132.960 1.120 ;
  LAYER metal4 ;
  RECT 1129.420 0.000 1132.960 1.120 ;
  LAYER metal3 ;
  RECT 1129.420 0.000 1132.960 1.120 ;
  LAYER metal2 ;
  RECT 1129.420 0.000 1132.960 1.120 ;
  LAYER metal1 ;
  RECT 1129.420 0.000 1132.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1115.780 0.000 1119.320 1.120 ;
  LAYER metal4 ;
  RECT 1115.780 0.000 1119.320 1.120 ;
  LAYER metal3 ;
  RECT 1115.780 0.000 1119.320 1.120 ;
  LAYER metal2 ;
  RECT 1115.780 0.000 1119.320 1.120 ;
  LAYER metal1 ;
  RECT 1115.780 0.000 1119.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1102.760 0.000 1106.300 1.120 ;
  LAYER metal4 ;
  RECT 1102.760 0.000 1106.300 1.120 ;
  LAYER metal3 ;
  RECT 1102.760 0.000 1106.300 1.120 ;
  LAYER metal2 ;
  RECT 1102.760 0.000 1106.300 1.120 ;
  LAYER metal1 ;
  RECT 1102.760 0.000 1106.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1035.180 0.000 1038.720 1.120 ;
  LAYER metal4 ;
  RECT 1035.180 0.000 1038.720 1.120 ;
  LAYER metal3 ;
  RECT 1035.180 0.000 1038.720 1.120 ;
  LAYER metal2 ;
  RECT 1035.180 0.000 1038.720 1.120 ;
  LAYER metal1 ;
  RECT 1035.180 0.000 1038.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1021.540 0.000 1025.080 1.120 ;
  LAYER metal4 ;
  RECT 1021.540 0.000 1025.080 1.120 ;
  LAYER metal3 ;
  RECT 1021.540 0.000 1025.080 1.120 ;
  LAYER metal2 ;
  RECT 1021.540 0.000 1025.080 1.120 ;
  LAYER metal1 ;
  RECT 1021.540 0.000 1025.080 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1010.380 0.000 1013.920 1.120 ;
  LAYER metal4 ;
  RECT 1010.380 0.000 1013.920 1.120 ;
  LAYER metal3 ;
  RECT 1010.380 0.000 1013.920 1.120 ;
  LAYER metal2 ;
  RECT 1010.380 0.000 1013.920 1.120 ;
  LAYER metal1 ;
  RECT 1010.380 0.000 1013.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 994.880 0.000 998.420 1.120 ;
  LAYER metal4 ;
  RECT 994.880 0.000 998.420 1.120 ;
  LAYER metal3 ;
  RECT 994.880 0.000 998.420 1.120 ;
  LAYER metal2 ;
  RECT 994.880 0.000 998.420 1.120 ;
  LAYER metal1 ;
  RECT 994.880 0.000 998.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 981.240 0.000 984.780 1.120 ;
  LAYER metal4 ;
  RECT 981.240 0.000 984.780 1.120 ;
  LAYER metal3 ;
  RECT 981.240 0.000 984.780 1.120 ;
  LAYER metal2 ;
  RECT 981.240 0.000 984.780 1.120 ;
  LAYER metal1 ;
  RECT 981.240 0.000 984.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 968.220 0.000 971.760 1.120 ;
  LAYER metal4 ;
  RECT 968.220 0.000 971.760 1.120 ;
  LAYER metal3 ;
  RECT 968.220 0.000 971.760 1.120 ;
  LAYER metal2 ;
  RECT 968.220 0.000 971.760 1.120 ;
  LAYER metal1 ;
  RECT 968.220 0.000 971.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 900.640 0.000 904.180 1.120 ;
  LAYER metal4 ;
  RECT 900.640 0.000 904.180 1.120 ;
  LAYER metal3 ;
  RECT 900.640 0.000 904.180 1.120 ;
  LAYER metal2 ;
  RECT 900.640 0.000 904.180 1.120 ;
  LAYER metal1 ;
  RECT 900.640 0.000 904.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 887.620 0.000 891.160 1.120 ;
  LAYER metal4 ;
  RECT 887.620 0.000 891.160 1.120 ;
  LAYER metal3 ;
  RECT 887.620 0.000 891.160 1.120 ;
  LAYER metal2 ;
  RECT 887.620 0.000 891.160 1.120 ;
  LAYER metal1 ;
  RECT 887.620 0.000 891.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 873.980 0.000 877.520 1.120 ;
  LAYER metal4 ;
  RECT 873.980 0.000 877.520 1.120 ;
  LAYER metal3 ;
  RECT 873.980 0.000 877.520 1.120 ;
  LAYER metal2 ;
  RECT 873.980 0.000 877.520 1.120 ;
  LAYER metal1 ;
  RECT 873.980 0.000 877.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 860.340 0.000 863.880 1.120 ;
  LAYER metal4 ;
  RECT 860.340 0.000 863.880 1.120 ;
  LAYER metal3 ;
  RECT 860.340 0.000 863.880 1.120 ;
  LAYER metal2 ;
  RECT 860.340 0.000 863.880 1.120 ;
  LAYER metal1 ;
  RECT 860.340 0.000 863.880 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 847.320 0.000 850.860 1.120 ;
  LAYER metal4 ;
  RECT 847.320 0.000 850.860 1.120 ;
  LAYER metal3 ;
  RECT 847.320 0.000 850.860 1.120 ;
  LAYER metal2 ;
  RECT 847.320 0.000 850.860 1.120 ;
  LAYER metal1 ;
  RECT 847.320 0.000 850.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 833.680 0.000 837.220 1.120 ;
  LAYER metal4 ;
  RECT 833.680 0.000 837.220 1.120 ;
  LAYER metal3 ;
  RECT 833.680 0.000 837.220 1.120 ;
  LAYER metal2 ;
  RECT 833.680 0.000 837.220 1.120 ;
  LAYER metal1 ;
  RECT 833.680 0.000 837.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 766.720 0.000 770.260 1.120 ;
  LAYER metal4 ;
  RECT 766.720 0.000 770.260 1.120 ;
  LAYER metal3 ;
  RECT 766.720 0.000 770.260 1.120 ;
  LAYER metal2 ;
  RECT 766.720 0.000 770.260 1.120 ;
  LAYER metal1 ;
  RECT 766.720 0.000 770.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 753.080 0.000 756.620 1.120 ;
  LAYER metal4 ;
  RECT 753.080 0.000 756.620 1.120 ;
  LAYER metal3 ;
  RECT 753.080 0.000 756.620 1.120 ;
  LAYER metal2 ;
  RECT 753.080 0.000 756.620 1.120 ;
  LAYER metal1 ;
  RECT 753.080 0.000 756.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 739.440 0.000 742.980 1.120 ;
  LAYER metal4 ;
  RECT 739.440 0.000 742.980 1.120 ;
  LAYER metal3 ;
  RECT 739.440 0.000 742.980 1.120 ;
  LAYER metal2 ;
  RECT 739.440 0.000 742.980 1.120 ;
  LAYER metal1 ;
  RECT 739.440 0.000 742.980 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 726.420 0.000 729.960 1.120 ;
  LAYER metal4 ;
  RECT 726.420 0.000 729.960 1.120 ;
  LAYER metal3 ;
  RECT 726.420 0.000 729.960 1.120 ;
  LAYER metal2 ;
  RECT 726.420 0.000 729.960 1.120 ;
  LAYER metal1 ;
  RECT 726.420 0.000 729.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 712.780 0.000 716.320 1.120 ;
  LAYER metal4 ;
  RECT 712.780 0.000 716.320 1.120 ;
  LAYER metal3 ;
  RECT 712.780 0.000 716.320 1.120 ;
  LAYER metal2 ;
  RECT 712.780 0.000 716.320 1.120 ;
  LAYER metal1 ;
  RECT 712.780 0.000 716.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 699.140 0.000 702.680 1.120 ;
  LAYER metal4 ;
  RECT 699.140 0.000 702.680 1.120 ;
  LAYER metal3 ;
  RECT 699.140 0.000 702.680 1.120 ;
  LAYER metal2 ;
  RECT 699.140 0.000 702.680 1.120 ;
  LAYER metal1 ;
  RECT 699.140 0.000 702.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 632.180 0.000 635.720 1.120 ;
  LAYER metal4 ;
  RECT 632.180 0.000 635.720 1.120 ;
  LAYER metal3 ;
  RECT 632.180 0.000 635.720 1.120 ;
  LAYER metal2 ;
  RECT 632.180 0.000 635.720 1.120 ;
  LAYER metal1 ;
  RECT 632.180 0.000 635.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 618.540 0.000 622.080 1.120 ;
  LAYER metal4 ;
  RECT 618.540 0.000 622.080 1.120 ;
  LAYER metal3 ;
  RECT 618.540 0.000 622.080 1.120 ;
  LAYER metal2 ;
  RECT 618.540 0.000 622.080 1.120 ;
  LAYER metal1 ;
  RECT 618.540 0.000 622.080 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 604.900 0.000 608.440 1.120 ;
  LAYER metal4 ;
  RECT 604.900 0.000 608.440 1.120 ;
  LAYER metal3 ;
  RECT 604.900 0.000 608.440 1.120 ;
  LAYER metal2 ;
  RECT 604.900 0.000 608.440 1.120 ;
  LAYER metal1 ;
  RECT 604.900 0.000 608.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 591.880 0.000 595.420 1.120 ;
  LAYER metal4 ;
  RECT 591.880 0.000 595.420 1.120 ;
  LAYER metal3 ;
  RECT 591.880 0.000 595.420 1.120 ;
  LAYER metal2 ;
  RECT 591.880 0.000 595.420 1.120 ;
  LAYER metal1 ;
  RECT 591.880 0.000 595.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 580.720 0.000 584.260 1.120 ;
  LAYER metal4 ;
  RECT 580.720 0.000 584.260 1.120 ;
  LAYER metal3 ;
  RECT 580.720 0.000 584.260 1.120 ;
  LAYER metal2 ;
  RECT 580.720 0.000 584.260 1.120 ;
  LAYER metal1 ;
  RECT 580.720 0.000 584.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 564.600 0.000 568.140 1.120 ;
  LAYER metal4 ;
  RECT 564.600 0.000 568.140 1.120 ;
  LAYER metal3 ;
  RECT 564.600 0.000 568.140 1.120 ;
  LAYER metal2 ;
  RECT 564.600 0.000 568.140 1.120 ;
  LAYER metal1 ;
  RECT 564.600 0.000 568.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 470.980 0.000 474.520 1.120 ;
  LAYER metal4 ;
  RECT 470.980 0.000 474.520 1.120 ;
  LAYER metal3 ;
  RECT 470.980 0.000 474.520 1.120 ;
  LAYER metal2 ;
  RECT 470.980 0.000 474.520 1.120 ;
  LAYER metal1 ;
  RECT 470.980 0.000 474.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 462.300 0.000 465.840 1.120 ;
  LAYER metal4 ;
  RECT 462.300 0.000 465.840 1.120 ;
  LAYER metal3 ;
  RECT 462.300 0.000 465.840 1.120 ;
  LAYER metal2 ;
  RECT 462.300 0.000 465.840 1.120 ;
  LAYER metal1 ;
  RECT 462.300 0.000 465.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 453.620 0.000 457.160 1.120 ;
  LAYER metal4 ;
  RECT 453.620 0.000 457.160 1.120 ;
  LAYER metal3 ;
  RECT 453.620 0.000 457.160 1.120 ;
  LAYER metal2 ;
  RECT 453.620 0.000 457.160 1.120 ;
  LAYER metal1 ;
  RECT 453.620 0.000 457.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 439.980 0.000 443.520 1.120 ;
  LAYER metal4 ;
  RECT 439.980 0.000 443.520 1.120 ;
  LAYER metal3 ;
  RECT 439.980 0.000 443.520 1.120 ;
  LAYER metal2 ;
  RECT 439.980 0.000 443.520 1.120 ;
  LAYER metal1 ;
  RECT 439.980 0.000 443.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER metal4 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER metal3 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER metal2 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER metal1 ;
  RECT 431.300 0.000 434.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 418.280 0.000 421.820 1.120 ;
  LAYER metal4 ;
  RECT 418.280 0.000 421.820 1.120 ;
  LAYER metal3 ;
  RECT 418.280 0.000 421.820 1.120 ;
  LAYER metal2 ;
  RECT 418.280 0.000 421.820 1.120 ;
  LAYER metal1 ;
  RECT 418.280 0.000 421.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 350.700 0.000 354.240 1.120 ;
  LAYER metal4 ;
  RECT 350.700 0.000 354.240 1.120 ;
  LAYER metal3 ;
  RECT 350.700 0.000 354.240 1.120 ;
  LAYER metal2 ;
  RECT 350.700 0.000 354.240 1.120 ;
  LAYER metal1 ;
  RECT 350.700 0.000 354.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 337.680 0.000 341.220 1.120 ;
  LAYER metal4 ;
  RECT 337.680 0.000 341.220 1.120 ;
  LAYER metal3 ;
  RECT 337.680 0.000 341.220 1.120 ;
  LAYER metal2 ;
  RECT 337.680 0.000 341.220 1.120 ;
  LAYER metal1 ;
  RECT 337.680 0.000 341.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 324.040 0.000 327.580 1.120 ;
  LAYER metal4 ;
  RECT 324.040 0.000 327.580 1.120 ;
  LAYER metal3 ;
  RECT 324.040 0.000 327.580 1.120 ;
  LAYER metal2 ;
  RECT 324.040 0.000 327.580 1.120 ;
  LAYER metal1 ;
  RECT 324.040 0.000 327.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 310.400 0.000 313.940 1.120 ;
  LAYER metal4 ;
  RECT 310.400 0.000 313.940 1.120 ;
  LAYER metal3 ;
  RECT 310.400 0.000 313.940 1.120 ;
  LAYER metal2 ;
  RECT 310.400 0.000 313.940 1.120 ;
  LAYER metal1 ;
  RECT 310.400 0.000 313.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 297.380 0.000 300.920 1.120 ;
  LAYER metal4 ;
  RECT 297.380 0.000 300.920 1.120 ;
  LAYER metal3 ;
  RECT 297.380 0.000 300.920 1.120 ;
  LAYER metal2 ;
  RECT 297.380 0.000 300.920 1.120 ;
  LAYER metal1 ;
  RECT 297.380 0.000 300.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 283.740 0.000 287.280 1.120 ;
  LAYER metal4 ;
  RECT 283.740 0.000 287.280 1.120 ;
  LAYER metal3 ;
  RECT 283.740 0.000 287.280 1.120 ;
  LAYER metal2 ;
  RECT 283.740 0.000 287.280 1.120 ;
  LAYER metal1 ;
  RECT 283.740 0.000 287.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 216.780 0.000 220.320 1.120 ;
  LAYER metal4 ;
  RECT 216.780 0.000 220.320 1.120 ;
  LAYER metal3 ;
  RECT 216.780 0.000 220.320 1.120 ;
  LAYER metal2 ;
  RECT 216.780 0.000 220.320 1.120 ;
  LAYER metal1 ;
  RECT 216.780 0.000 220.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 203.140 0.000 206.680 1.120 ;
  LAYER metal4 ;
  RECT 203.140 0.000 206.680 1.120 ;
  LAYER metal3 ;
  RECT 203.140 0.000 206.680 1.120 ;
  LAYER metal2 ;
  RECT 203.140 0.000 206.680 1.120 ;
  LAYER metal1 ;
  RECT 203.140 0.000 206.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 189.500 0.000 193.040 1.120 ;
  LAYER metal4 ;
  RECT 189.500 0.000 193.040 1.120 ;
  LAYER metal3 ;
  RECT 189.500 0.000 193.040 1.120 ;
  LAYER metal2 ;
  RECT 189.500 0.000 193.040 1.120 ;
  LAYER metal1 ;
  RECT 189.500 0.000 193.040 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER metal4 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER metal3 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER metal2 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER metal1 ;
  RECT 176.480 0.000 180.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 162.840 0.000 166.380 1.120 ;
  LAYER metal4 ;
  RECT 162.840 0.000 166.380 1.120 ;
  LAYER metal3 ;
  RECT 162.840 0.000 166.380 1.120 ;
  LAYER metal2 ;
  RECT 162.840 0.000 166.380 1.120 ;
  LAYER metal1 ;
  RECT 162.840 0.000 166.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 149.200 0.000 152.740 1.120 ;
  LAYER metal4 ;
  RECT 149.200 0.000 152.740 1.120 ;
  LAYER metal3 ;
  RECT 149.200 0.000 152.740 1.120 ;
  LAYER metal2 ;
  RECT 149.200 0.000 152.740 1.120 ;
  LAYER metal1 ;
  RECT 149.200 0.000 152.740 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 82.240 0.000 85.780 1.120 ;
  LAYER metal4 ;
  RECT 82.240 0.000 85.780 1.120 ;
  LAYER metal3 ;
  RECT 82.240 0.000 85.780 1.120 ;
  LAYER metal2 ;
  RECT 82.240 0.000 85.780 1.120 ;
  LAYER metal1 ;
  RECT 82.240 0.000 85.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 68.600 0.000 72.140 1.120 ;
  LAYER metal4 ;
  RECT 68.600 0.000 72.140 1.120 ;
  LAYER metal3 ;
  RECT 68.600 0.000 72.140 1.120 ;
  LAYER metal2 ;
  RECT 68.600 0.000 72.140 1.120 ;
  LAYER metal1 ;
  RECT 68.600 0.000 72.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER metal4 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER metal3 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER metal2 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER metal1 ;
  RECT 54.960 0.000 58.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER metal4 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER metal3 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER metal2 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER metal1 ;
  RECT 41.940 0.000 45.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER metal4 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER metal3 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER metal2 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER metal1 ;
  RECT 28.300 0.000 31.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 17.140 0.000 20.680 1.120 ;
  LAYER metal4 ;
  RECT 17.140 0.000 20.680 1.120 ;
  LAYER metal3 ;
  RECT 17.140 0.000 20.680 1.120 ;
  LAYER metal2 ;
  RECT 17.140 0.000 20.680 1.120 ;
  LAYER metal1 ;
  RECT 17.140 0.000 20.680 1.120 ;
 END
END GND
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal5 ;
  RECT 1444.720 517.220 1445.840 520.460 ;
  LAYER metal4 ;
  RECT 1444.720 517.220 1445.840 520.460 ;
  LAYER metal3 ;
  RECT 1444.720 517.220 1445.840 520.460 ;
  LAYER metal2 ;
  RECT 1444.720 517.220 1445.840 520.460 ;
  LAYER metal1 ;
  RECT 1444.720 517.220 1445.840 520.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 509.380 1445.840 512.620 ;
  LAYER metal4 ;
  RECT 1444.720 509.380 1445.840 512.620 ;
  LAYER metal3 ;
  RECT 1444.720 509.380 1445.840 512.620 ;
  LAYER metal2 ;
  RECT 1444.720 509.380 1445.840 512.620 ;
  LAYER metal1 ;
  RECT 1444.720 509.380 1445.840 512.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 501.540 1445.840 504.780 ;
  LAYER metal4 ;
  RECT 1444.720 501.540 1445.840 504.780 ;
  LAYER metal3 ;
  RECT 1444.720 501.540 1445.840 504.780 ;
  LAYER metal2 ;
  RECT 1444.720 501.540 1445.840 504.780 ;
  LAYER metal1 ;
  RECT 1444.720 501.540 1445.840 504.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 493.700 1445.840 496.940 ;
  LAYER metal4 ;
  RECT 1444.720 493.700 1445.840 496.940 ;
  LAYER metal3 ;
  RECT 1444.720 493.700 1445.840 496.940 ;
  LAYER metal2 ;
  RECT 1444.720 493.700 1445.840 496.940 ;
  LAYER metal1 ;
  RECT 1444.720 493.700 1445.840 496.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 485.860 1445.840 489.100 ;
  LAYER metal4 ;
  RECT 1444.720 485.860 1445.840 489.100 ;
  LAYER metal3 ;
  RECT 1444.720 485.860 1445.840 489.100 ;
  LAYER metal2 ;
  RECT 1444.720 485.860 1445.840 489.100 ;
  LAYER metal1 ;
  RECT 1444.720 485.860 1445.840 489.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 478.020 1445.840 481.260 ;
  LAYER metal4 ;
  RECT 1444.720 478.020 1445.840 481.260 ;
  LAYER metal3 ;
  RECT 1444.720 478.020 1445.840 481.260 ;
  LAYER metal2 ;
  RECT 1444.720 478.020 1445.840 481.260 ;
  LAYER metal1 ;
  RECT 1444.720 478.020 1445.840 481.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 438.820 1445.840 442.060 ;
  LAYER metal4 ;
  RECT 1444.720 438.820 1445.840 442.060 ;
  LAYER metal3 ;
  RECT 1444.720 438.820 1445.840 442.060 ;
  LAYER metal2 ;
  RECT 1444.720 438.820 1445.840 442.060 ;
  LAYER metal1 ;
  RECT 1444.720 438.820 1445.840 442.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 430.980 1445.840 434.220 ;
  LAYER metal4 ;
  RECT 1444.720 430.980 1445.840 434.220 ;
  LAYER metal3 ;
  RECT 1444.720 430.980 1445.840 434.220 ;
  LAYER metal2 ;
  RECT 1444.720 430.980 1445.840 434.220 ;
  LAYER metal1 ;
  RECT 1444.720 430.980 1445.840 434.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 423.140 1445.840 426.380 ;
  LAYER metal4 ;
  RECT 1444.720 423.140 1445.840 426.380 ;
  LAYER metal3 ;
  RECT 1444.720 423.140 1445.840 426.380 ;
  LAYER metal2 ;
  RECT 1444.720 423.140 1445.840 426.380 ;
  LAYER metal1 ;
  RECT 1444.720 423.140 1445.840 426.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 415.300 1445.840 418.540 ;
  LAYER metal4 ;
  RECT 1444.720 415.300 1445.840 418.540 ;
  LAYER metal3 ;
  RECT 1444.720 415.300 1445.840 418.540 ;
  LAYER metal2 ;
  RECT 1444.720 415.300 1445.840 418.540 ;
  LAYER metal1 ;
  RECT 1444.720 415.300 1445.840 418.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 407.460 1445.840 410.700 ;
  LAYER metal4 ;
  RECT 1444.720 407.460 1445.840 410.700 ;
  LAYER metal3 ;
  RECT 1444.720 407.460 1445.840 410.700 ;
  LAYER metal2 ;
  RECT 1444.720 407.460 1445.840 410.700 ;
  LAYER metal1 ;
  RECT 1444.720 407.460 1445.840 410.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 399.620 1445.840 402.860 ;
  LAYER metal4 ;
  RECT 1444.720 399.620 1445.840 402.860 ;
  LAYER metal3 ;
  RECT 1444.720 399.620 1445.840 402.860 ;
  LAYER metal2 ;
  RECT 1444.720 399.620 1445.840 402.860 ;
  LAYER metal1 ;
  RECT 1444.720 399.620 1445.840 402.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 360.420 1445.840 363.660 ;
  LAYER metal4 ;
  RECT 1444.720 360.420 1445.840 363.660 ;
  LAYER metal3 ;
  RECT 1444.720 360.420 1445.840 363.660 ;
  LAYER metal2 ;
  RECT 1444.720 360.420 1445.840 363.660 ;
  LAYER metal1 ;
  RECT 1444.720 360.420 1445.840 363.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 352.580 1445.840 355.820 ;
  LAYER metal4 ;
  RECT 1444.720 352.580 1445.840 355.820 ;
  LAYER metal3 ;
  RECT 1444.720 352.580 1445.840 355.820 ;
  LAYER metal2 ;
  RECT 1444.720 352.580 1445.840 355.820 ;
  LAYER metal1 ;
  RECT 1444.720 352.580 1445.840 355.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 344.740 1445.840 347.980 ;
  LAYER metal4 ;
  RECT 1444.720 344.740 1445.840 347.980 ;
  LAYER metal3 ;
  RECT 1444.720 344.740 1445.840 347.980 ;
  LAYER metal2 ;
  RECT 1444.720 344.740 1445.840 347.980 ;
  LAYER metal1 ;
  RECT 1444.720 344.740 1445.840 347.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 336.900 1445.840 340.140 ;
  LAYER metal4 ;
  RECT 1444.720 336.900 1445.840 340.140 ;
  LAYER metal3 ;
  RECT 1444.720 336.900 1445.840 340.140 ;
  LAYER metal2 ;
  RECT 1444.720 336.900 1445.840 340.140 ;
  LAYER metal1 ;
  RECT 1444.720 336.900 1445.840 340.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 329.060 1445.840 332.300 ;
  LAYER metal4 ;
  RECT 1444.720 329.060 1445.840 332.300 ;
  LAYER metal3 ;
  RECT 1444.720 329.060 1445.840 332.300 ;
  LAYER metal2 ;
  RECT 1444.720 329.060 1445.840 332.300 ;
  LAYER metal1 ;
  RECT 1444.720 329.060 1445.840 332.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 321.220 1445.840 324.460 ;
  LAYER metal4 ;
  RECT 1444.720 321.220 1445.840 324.460 ;
  LAYER metal3 ;
  RECT 1444.720 321.220 1445.840 324.460 ;
  LAYER metal2 ;
  RECT 1444.720 321.220 1445.840 324.460 ;
  LAYER metal1 ;
  RECT 1444.720 321.220 1445.840 324.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 282.020 1445.840 285.260 ;
  LAYER metal4 ;
  RECT 1444.720 282.020 1445.840 285.260 ;
  LAYER metal3 ;
  RECT 1444.720 282.020 1445.840 285.260 ;
  LAYER metal2 ;
  RECT 1444.720 282.020 1445.840 285.260 ;
  LAYER metal1 ;
  RECT 1444.720 282.020 1445.840 285.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 274.180 1445.840 277.420 ;
  LAYER metal4 ;
  RECT 1444.720 274.180 1445.840 277.420 ;
  LAYER metal3 ;
  RECT 1444.720 274.180 1445.840 277.420 ;
  LAYER metal2 ;
  RECT 1444.720 274.180 1445.840 277.420 ;
  LAYER metal1 ;
  RECT 1444.720 274.180 1445.840 277.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 266.340 1445.840 269.580 ;
  LAYER metal4 ;
  RECT 1444.720 266.340 1445.840 269.580 ;
  LAYER metal3 ;
  RECT 1444.720 266.340 1445.840 269.580 ;
  LAYER metal2 ;
  RECT 1444.720 266.340 1445.840 269.580 ;
  LAYER metal1 ;
  RECT 1444.720 266.340 1445.840 269.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 258.500 1445.840 261.740 ;
  LAYER metal4 ;
  RECT 1444.720 258.500 1445.840 261.740 ;
  LAYER metal3 ;
  RECT 1444.720 258.500 1445.840 261.740 ;
  LAYER metal2 ;
  RECT 1444.720 258.500 1445.840 261.740 ;
  LAYER metal1 ;
  RECT 1444.720 258.500 1445.840 261.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 250.660 1445.840 253.900 ;
  LAYER metal4 ;
  RECT 1444.720 250.660 1445.840 253.900 ;
  LAYER metal3 ;
  RECT 1444.720 250.660 1445.840 253.900 ;
  LAYER metal2 ;
  RECT 1444.720 250.660 1445.840 253.900 ;
  LAYER metal1 ;
  RECT 1444.720 250.660 1445.840 253.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 242.820 1445.840 246.060 ;
  LAYER metal4 ;
  RECT 1444.720 242.820 1445.840 246.060 ;
  LAYER metal3 ;
  RECT 1444.720 242.820 1445.840 246.060 ;
  LAYER metal2 ;
  RECT 1444.720 242.820 1445.840 246.060 ;
  LAYER metal1 ;
  RECT 1444.720 242.820 1445.840 246.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 203.620 1445.840 206.860 ;
  LAYER metal4 ;
  RECT 1444.720 203.620 1445.840 206.860 ;
  LAYER metal3 ;
  RECT 1444.720 203.620 1445.840 206.860 ;
  LAYER metal2 ;
  RECT 1444.720 203.620 1445.840 206.860 ;
  LAYER metal1 ;
  RECT 1444.720 203.620 1445.840 206.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 195.780 1445.840 199.020 ;
  LAYER metal4 ;
  RECT 1444.720 195.780 1445.840 199.020 ;
  LAYER metal3 ;
  RECT 1444.720 195.780 1445.840 199.020 ;
  LAYER metal2 ;
  RECT 1444.720 195.780 1445.840 199.020 ;
  LAYER metal1 ;
  RECT 1444.720 195.780 1445.840 199.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 187.940 1445.840 191.180 ;
  LAYER metal4 ;
  RECT 1444.720 187.940 1445.840 191.180 ;
  LAYER metal3 ;
  RECT 1444.720 187.940 1445.840 191.180 ;
  LAYER metal2 ;
  RECT 1444.720 187.940 1445.840 191.180 ;
  LAYER metal1 ;
  RECT 1444.720 187.940 1445.840 191.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 180.100 1445.840 183.340 ;
  LAYER metal4 ;
  RECT 1444.720 180.100 1445.840 183.340 ;
  LAYER metal3 ;
  RECT 1444.720 180.100 1445.840 183.340 ;
  LAYER metal2 ;
  RECT 1444.720 180.100 1445.840 183.340 ;
  LAYER metal1 ;
  RECT 1444.720 180.100 1445.840 183.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 172.260 1445.840 175.500 ;
  LAYER metal4 ;
  RECT 1444.720 172.260 1445.840 175.500 ;
  LAYER metal3 ;
  RECT 1444.720 172.260 1445.840 175.500 ;
  LAYER metal2 ;
  RECT 1444.720 172.260 1445.840 175.500 ;
  LAYER metal1 ;
  RECT 1444.720 172.260 1445.840 175.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 164.420 1445.840 167.660 ;
  LAYER metal4 ;
  RECT 1444.720 164.420 1445.840 167.660 ;
  LAYER metal3 ;
  RECT 1444.720 164.420 1445.840 167.660 ;
  LAYER metal2 ;
  RECT 1444.720 164.420 1445.840 167.660 ;
  LAYER metal1 ;
  RECT 1444.720 164.420 1445.840 167.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 125.220 1445.840 128.460 ;
  LAYER metal4 ;
  RECT 1444.720 125.220 1445.840 128.460 ;
  LAYER metal3 ;
  RECT 1444.720 125.220 1445.840 128.460 ;
  LAYER metal2 ;
  RECT 1444.720 125.220 1445.840 128.460 ;
  LAYER metal1 ;
  RECT 1444.720 125.220 1445.840 128.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 117.380 1445.840 120.620 ;
  LAYER metal4 ;
  RECT 1444.720 117.380 1445.840 120.620 ;
  LAYER metal3 ;
  RECT 1444.720 117.380 1445.840 120.620 ;
  LAYER metal2 ;
  RECT 1444.720 117.380 1445.840 120.620 ;
  LAYER metal1 ;
  RECT 1444.720 117.380 1445.840 120.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 109.540 1445.840 112.780 ;
  LAYER metal4 ;
  RECT 1444.720 109.540 1445.840 112.780 ;
  LAYER metal3 ;
  RECT 1444.720 109.540 1445.840 112.780 ;
  LAYER metal2 ;
  RECT 1444.720 109.540 1445.840 112.780 ;
  LAYER metal1 ;
  RECT 1444.720 109.540 1445.840 112.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 101.700 1445.840 104.940 ;
  LAYER metal4 ;
  RECT 1444.720 101.700 1445.840 104.940 ;
  LAYER metal3 ;
  RECT 1444.720 101.700 1445.840 104.940 ;
  LAYER metal2 ;
  RECT 1444.720 101.700 1445.840 104.940 ;
  LAYER metal1 ;
  RECT 1444.720 101.700 1445.840 104.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 93.860 1445.840 97.100 ;
  LAYER metal4 ;
  RECT 1444.720 93.860 1445.840 97.100 ;
  LAYER metal3 ;
  RECT 1444.720 93.860 1445.840 97.100 ;
  LAYER metal2 ;
  RECT 1444.720 93.860 1445.840 97.100 ;
  LAYER metal1 ;
  RECT 1444.720 93.860 1445.840 97.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 86.020 1445.840 89.260 ;
  LAYER metal4 ;
  RECT 1444.720 86.020 1445.840 89.260 ;
  LAYER metal3 ;
  RECT 1444.720 86.020 1445.840 89.260 ;
  LAYER metal2 ;
  RECT 1444.720 86.020 1445.840 89.260 ;
  LAYER metal1 ;
  RECT 1444.720 86.020 1445.840 89.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 46.820 1445.840 50.060 ;
  LAYER metal4 ;
  RECT 1444.720 46.820 1445.840 50.060 ;
  LAYER metal3 ;
  RECT 1444.720 46.820 1445.840 50.060 ;
  LAYER metal2 ;
  RECT 1444.720 46.820 1445.840 50.060 ;
  LAYER metal1 ;
  RECT 1444.720 46.820 1445.840 50.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 38.980 1445.840 42.220 ;
  LAYER metal4 ;
  RECT 1444.720 38.980 1445.840 42.220 ;
  LAYER metal3 ;
  RECT 1444.720 38.980 1445.840 42.220 ;
  LAYER metal2 ;
  RECT 1444.720 38.980 1445.840 42.220 ;
  LAYER metal1 ;
  RECT 1444.720 38.980 1445.840 42.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 31.140 1445.840 34.380 ;
  LAYER metal4 ;
  RECT 1444.720 31.140 1445.840 34.380 ;
  LAYER metal3 ;
  RECT 1444.720 31.140 1445.840 34.380 ;
  LAYER metal2 ;
  RECT 1444.720 31.140 1445.840 34.380 ;
  LAYER metal1 ;
  RECT 1444.720 31.140 1445.840 34.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 23.300 1445.840 26.540 ;
  LAYER metal4 ;
  RECT 1444.720 23.300 1445.840 26.540 ;
  LAYER metal3 ;
  RECT 1444.720 23.300 1445.840 26.540 ;
  LAYER metal2 ;
  RECT 1444.720 23.300 1445.840 26.540 ;
  LAYER metal1 ;
  RECT 1444.720 23.300 1445.840 26.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 15.460 1445.840 18.700 ;
  LAYER metal4 ;
  RECT 1444.720 15.460 1445.840 18.700 ;
  LAYER metal3 ;
  RECT 1444.720 15.460 1445.840 18.700 ;
  LAYER metal2 ;
  RECT 1444.720 15.460 1445.840 18.700 ;
  LAYER metal1 ;
  RECT 1444.720 15.460 1445.840 18.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1444.720 7.620 1445.840 10.860 ;
  LAYER metal4 ;
  RECT 1444.720 7.620 1445.840 10.860 ;
  LAYER metal3 ;
  RECT 1444.720 7.620 1445.840 10.860 ;
  LAYER metal2 ;
  RECT 1444.720 7.620 1445.840 10.860 ;
  LAYER metal1 ;
  RECT 1444.720 7.620 1445.840 10.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 517.220 1.120 520.460 ;
  LAYER metal4 ;
  RECT 0.000 517.220 1.120 520.460 ;
  LAYER metal3 ;
  RECT 0.000 517.220 1.120 520.460 ;
  LAYER metal2 ;
  RECT 0.000 517.220 1.120 520.460 ;
  LAYER metal1 ;
  RECT 0.000 517.220 1.120 520.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 509.380 1.120 512.620 ;
  LAYER metal4 ;
  RECT 0.000 509.380 1.120 512.620 ;
  LAYER metal3 ;
  RECT 0.000 509.380 1.120 512.620 ;
  LAYER metal2 ;
  RECT 0.000 509.380 1.120 512.620 ;
  LAYER metal1 ;
  RECT 0.000 509.380 1.120 512.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 501.540 1.120 504.780 ;
  LAYER metal4 ;
  RECT 0.000 501.540 1.120 504.780 ;
  LAYER metal3 ;
  RECT 0.000 501.540 1.120 504.780 ;
  LAYER metal2 ;
  RECT 0.000 501.540 1.120 504.780 ;
  LAYER metal1 ;
  RECT 0.000 501.540 1.120 504.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 493.700 1.120 496.940 ;
  LAYER metal4 ;
  RECT 0.000 493.700 1.120 496.940 ;
  LAYER metal3 ;
  RECT 0.000 493.700 1.120 496.940 ;
  LAYER metal2 ;
  RECT 0.000 493.700 1.120 496.940 ;
  LAYER metal1 ;
  RECT 0.000 493.700 1.120 496.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 485.860 1.120 489.100 ;
  LAYER metal4 ;
  RECT 0.000 485.860 1.120 489.100 ;
  LAYER metal3 ;
  RECT 0.000 485.860 1.120 489.100 ;
  LAYER metal2 ;
  RECT 0.000 485.860 1.120 489.100 ;
  LAYER metal1 ;
  RECT 0.000 485.860 1.120 489.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 478.020 1.120 481.260 ;
  LAYER metal4 ;
  RECT 0.000 478.020 1.120 481.260 ;
  LAYER metal3 ;
  RECT 0.000 478.020 1.120 481.260 ;
  LAYER metal2 ;
  RECT 0.000 478.020 1.120 481.260 ;
  LAYER metal1 ;
  RECT 0.000 478.020 1.120 481.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 438.820 1.120 442.060 ;
  LAYER metal4 ;
  RECT 0.000 438.820 1.120 442.060 ;
  LAYER metal3 ;
  RECT 0.000 438.820 1.120 442.060 ;
  LAYER metal2 ;
  RECT 0.000 438.820 1.120 442.060 ;
  LAYER metal1 ;
  RECT 0.000 438.820 1.120 442.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 430.980 1.120 434.220 ;
  LAYER metal4 ;
  RECT 0.000 430.980 1.120 434.220 ;
  LAYER metal3 ;
  RECT 0.000 430.980 1.120 434.220 ;
  LAYER metal2 ;
  RECT 0.000 430.980 1.120 434.220 ;
  LAYER metal1 ;
  RECT 0.000 430.980 1.120 434.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 423.140 1.120 426.380 ;
  LAYER metal4 ;
  RECT 0.000 423.140 1.120 426.380 ;
  LAYER metal3 ;
  RECT 0.000 423.140 1.120 426.380 ;
  LAYER metal2 ;
  RECT 0.000 423.140 1.120 426.380 ;
  LAYER metal1 ;
  RECT 0.000 423.140 1.120 426.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 415.300 1.120 418.540 ;
  LAYER metal4 ;
  RECT 0.000 415.300 1.120 418.540 ;
  LAYER metal3 ;
  RECT 0.000 415.300 1.120 418.540 ;
  LAYER metal2 ;
  RECT 0.000 415.300 1.120 418.540 ;
  LAYER metal1 ;
  RECT 0.000 415.300 1.120 418.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 407.460 1.120 410.700 ;
  LAYER metal4 ;
  RECT 0.000 407.460 1.120 410.700 ;
  LAYER metal3 ;
  RECT 0.000 407.460 1.120 410.700 ;
  LAYER metal2 ;
  RECT 0.000 407.460 1.120 410.700 ;
  LAYER metal1 ;
  RECT 0.000 407.460 1.120 410.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 399.620 1.120 402.860 ;
  LAYER metal4 ;
  RECT 0.000 399.620 1.120 402.860 ;
  LAYER metal3 ;
  RECT 0.000 399.620 1.120 402.860 ;
  LAYER metal2 ;
  RECT 0.000 399.620 1.120 402.860 ;
  LAYER metal1 ;
  RECT 0.000 399.620 1.120 402.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 360.420 1.120 363.660 ;
  LAYER metal4 ;
  RECT 0.000 360.420 1.120 363.660 ;
  LAYER metal3 ;
  RECT 0.000 360.420 1.120 363.660 ;
  LAYER metal2 ;
  RECT 0.000 360.420 1.120 363.660 ;
  LAYER metal1 ;
  RECT 0.000 360.420 1.120 363.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 352.580 1.120 355.820 ;
  LAYER metal4 ;
  RECT 0.000 352.580 1.120 355.820 ;
  LAYER metal3 ;
  RECT 0.000 352.580 1.120 355.820 ;
  LAYER metal2 ;
  RECT 0.000 352.580 1.120 355.820 ;
  LAYER metal1 ;
  RECT 0.000 352.580 1.120 355.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 344.740 1.120 347.980 ;
  LAYER metal4 ;
  RECT 0.000 344.740 1.120 347.980 ;
  LAYER metal3 ;
  RECT 0.000 344.740 1.120 347.980 ;
  LAYER metal2 ;
  RECT 0.000 344.740 1.120 347.980 ;
  LAYER metal1 ;
  RECT 0.000 344.740 1.120 347.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 336.900 1.120 340.140 ;
  LAYER metal4 ;
  RECT 0.000 336.900 1.120 340.140 ;
  LAYER metal3 ;
  RECT 0.000 336.900 1.120 340.140 ;
  LAYER metal2 ;
  RECT 0.000 336.900 1.120 340.140 ;
  LAYER metal1 ;
  RECT 0.000 336.900 1.120 340.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 329.060 1.120 332.300 ;
  LAYER metal4 ;
  RECT 0.000 329.060 1.120 332.300 ;
  LAYER metal3 ;
  RECT 0.000 329.060 1.120 332.300 ;
  LAYER metal2 ;
  RECT 0.000 329.060 1.120 332.300 ;
  LAYER metal1 ;
  RECT 0.000 329.060 1.120 332.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 321.220 1.120 324.460 ;
  LAYER metal4 ;
  RECT 0.000 321.220 1.120 324.460 ;
  LAYER metal3 ;
  RECT 0.000 321.220 1.120 324.460 ;
  LAYER metal2 ;
  RECT 0.000 321.220 1.120 324.460 ;
  LAYER metal1 ;
  RECT 0.000 321.220 1.120 324.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 282.020 1.120 285.260 ;
  LAYER metal4 ;
  RECT 0.000 282.020 1.120 285.260 ;
  LAYER metal3 ;
  RECT 0.000 282.020 1.120 285.260 ;
  LAYER metal2 ;
  RECT 0.000 282.020 1.120 285.260 ;
  LAYER metal1 ;
  RECT 0.000 282.020 1.120 285.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 274.180 1.120 277.420 ;
  LAYER metal4 ;
  RECT 0.000 274.180 1.120 277.420 ;
  LAYER metal3 ;
  RECT 0.000 274.180 1.120 277.420 ;
  LAYER metal2 ;
  RECT 0.000 274.180 1.120 277.420 ;
  LAYER metal1 ;
  RECT 0.000 274.180 1.120 277.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 266.340 1.120 269.580 ;
  LAYER metal4 ;
  RECT 0.000 266.340 1.120 269.580 ;
  LAYER metal3 ;
  RECT 0.000 266.340 1.120 269.580 ;
  LAYER metal2 ;
  RECT 0.000 266.340 1.120 269.580 ;
  LAYER metal1 ;
  RECT 0.000 266.340 1.120 269.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 258.500 1.120 261.740 ;
  LAYER metal4 ;
  RECT 0.000 258.500 1.120 261.740 ;
  LAYER metal3 ;
  RECT 0.000 258.500 1.120 261.740 ;
  LAYER metal2 ;
  RECT 0.000 258.500 1.120 261.740 ;
  LAYER metal1 ;
  RECT 0.000 258.500 1.120 261.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 250.660 1.120 253.900 ;
  LAYER metal4 ;
  RECT 0.000 250.660 1.120 253.900 ;
  LAYER metal3 ;
  RECT 0.000 250.660 1.120 253.900 ;
  LAYER metal2 ;
  RECT 0.000 250.660 1.120 253.900 ;
  LAYER metal1 ;
  RECT 0.000 250.660 1.120 253.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 242.820 1.120 246.060 ;
  LAYER metal4 ;
  RECT 0.000 242.820 1.120 246.060 ;
  LAYER metal3 ;
  RECT 0.000 242.820 1.120 246.060 ;
  LAYER metal2 ;
  RECT 0.000 242.820 1.120 246.060 ;
  LAYER metal1 ;
  RECT 0.000 242.820 1.120 246.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 203.620 1.120 206.860 ;
  LAYER metal4 ;
  RECT 0.000 203.620 1.120 206.860 ;
  LAYER metal3 ;
  RECT 0.000 203.620 1.120 206.860 ;
  LAYER metal2 ;
  RECT 0.000 203.620 1.120 206.860 ;
  LAYER metal1 ;
  RECT 0.000 203.620 1.120 206.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER metal4 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER metal3 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER metal2 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER metal1 ;
  RECT 0.000 195.780 1.120 199.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER metal4 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER metal3 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER metal2 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER metal1 ;
  RECT 0.000 187.940 1.120 191.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER metal4 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER metal3 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER metal2 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER metal1 ;
  RECT 0.000 180.100 1.120 183.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER metal4 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER metal3 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER metal2 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER metal1 ;
  RECT 0.000 172.260 1.120 175.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER metal4 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER metal3 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER metal2 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER metal1 ;
  RECT 0.000 164.420 1.120 167.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER metal4 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER metal3 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER metal2 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER metal1 ;
  RECT 0.000 125.220 1.120 128.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER metal4 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER metal3 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER metal2 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER metal1 ;
  RECT 0.000 117.380 1.120 120.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER metal4 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER metal3 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER metal2 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER metal1 ;
  RECT 0.000 109.540 1.120 112.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER metal4 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER metal3 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER metal2 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER metal1 ;
  RECT 0.000 101.700 1.120 104.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER metal4 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER metal3 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER metal2 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER metal1 ;
  RECT 0.000 93.860 1.120 97.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER metal4 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER metal3 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER metal2 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER metal1 ;
  RECT 0.000 86.020 1.120 89.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER metal4 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER metal3 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER metal2 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER metal1 ;
  RECT 0.000 46.820 1.120 50.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER metal4 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER metal3 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER metal2 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER metal1 ;
  RECT 0.000 38.980 1.120 42.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER metal4 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER metal3 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER metal2 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER metal1 ;
  RECT 0.000 31.140 1.120 34.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER metal4 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER metal3 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER metal2 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER metal1 ;
  RECT 0.000 23.300 1.120 26.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER metal4 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER metal3 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER metal2 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER metal1 ;
  RECT 0.000 15.460 1.120 18.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER metal4 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER metal3 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER metal2 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER metal1 ;
  RECT 0.000 7.620 1.120 10.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1429.500 543.200 1433.040 544.320 ;
  LAYER metal4 ;
  RECT 1429.500 543.200 1433.040 544.320 ;
  LAYER metal3 ;
  RECT 1429.500 543.200 1433.040 544.320 ;
  LAYER metal2 ;
  RECT 1429.500 543.200 1433.040 544.320 ;
  LAYER metal1 ;
  RECT 1429.500 543.200 1433.040 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1415.860 543.200 1419.400 544.320 ;
  LAYER metal4 ;
  RECT 1415.860 543.200 1419.400 544.320 ;
  LAYER metal3 ;
  RECT 1415.860 543.200 1419.400 544.320 ;
  LAYER metal2 ;
  RECT 1415.860 543.200 1419.400 544.320 ;
  LAYER metal1 ;
  RECT 1415.860 543.200 1419.400 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1402.220 543.200 1405.760 544.320 ;
  LAYER metal4 ;
  RECT 1402.220 543.200 1405.760 544.320 ;
  LAYER metal3 ;
  RECT 1402.220 543.200 1405.760 544.320 ;
  LAYER metal2 ;
  RECT 1402.220 543.200 1405.760 544.320 ;
  LAYER metal1 ;
  RECT 1402.220 543.200 1405.760 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1389.200 543.200 1392.740 544.320 ;
  LAYER metal4 ;
  RECT 1389.200 543.200 1392.740 544.320 ;
  LAYER metal3 ;
  RECT 1389.200 543.200 1392.740 544.320 ;
  LAYER metal2 ;
  RECT 1389.200 543.200 1392.740 544.320 ;
  LAYER metal1 ;
  RECT 1389.200 543.200 1392.740 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1375.560 543.200 1379.100 544.320 ;
  LAYER metal4 ;
  RECT 1375.560 543.200 1379.100 544.320 ;
  LAYER metal3 ;
  RECT 1375.560 543.200 1379.100 544.320 ;
  LAYER metal2 ;
  RECT 1375.560 543.200 1379.100 544.320 ;
  LAYER metal1 ;
  RECT 1375.560 543.200 1379.100 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1361.920 543.200 1365.460 544.320 ;
  LAYER metal4 ;
  RECT 1361.920 543.200 1365.460 544.320 ;
  LAYER metal3 ;
  RECT 1361.920 543.200 1365.460 544.320 ;
  LAYER metal2 ;
  RECT 1361.920 543.200 1365.460 544.320 ;
  LAYER metal1 ;
  RECT 1361.920 543.200 1365.460 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1294.960 543.200 1298.500 544.320 ;
  LAYER metal4 ;
  RECT 1294.960 543.200 1298.500 544.320 ;
  LAYER metal3 ;
  RECT 1294.960 543.200 1298.500 544.320 ;
  LAYER metal2 ;
  RECT 1294.960 543.200 1298.500 544.320 ;
  LAYER metal1 ;
  RECT 1294.960 543.200 1298.500 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1281.320 543.200 1284.860 544.320 ;
  LAYER metal4 ;
  RECT 1281.320 543.200 1284.860 544.320 ;
  LAYER metal3 ;
  RECT 1281.320 543.200 1284.860 544.320 ;
  LAYER metal2 ;
  RECT 1281.320 543.200 1284.860 544.320 ;
  LAYER metal1 ;
  RECT 1281.320 543.200 1284.860 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1268.300 543.200 1271.840 544.320 ;
  LAYER metal4 ;
  RECT 1268.300 543.200 1271.840 544.320 ;
  LAYER metal3 ;
  RECT 1268.300 543.200 1271.840 544.320 ;
  LAYER metal2 ;
  RECT 1268.300 543.200 1271.840 544.320 ;
  LAYER metal1 ;
  RECT 1268.300 543.200 1271.840 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1254.660 543.200 1258.200 544.320 ;
  LAYER metal4 ;
  RECT 1254.660 543.200 1258.200 544.320 ;
  LAYER metal3 ;
  RECT 1254.660 543.200 1258.200 544.320 ;
  LAYER metal2 ;
  RECT 1254.660 543.200 1258.200 544.320 ;
  LAYER metal1 ;
  RECT 1254.660 543.200 1258.200 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1241.020 543.200 1244.560 544.320 ;
  LAYER metal4 ;
  RECT 1241.020 543.200 1244.560 544.320 ;
  LAYER metal3 ;
  RECT 1241.020 543.200 1244.560 544.320 ;
  LAYER metal2 ;
  RECT 1241.020 543.200 1244.560 544.320 ;
  LAYER metal1 ;
  RECT 1241.020 543.200 1244.560 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1228.000 543.200 1231.540 544.320 ;
  LAYER metal4 ;
  RECT 1228.000 543.200 1231.540 544.320 ;
  LAYER metal3 ;
  RECT 1228.000 543.200 1231.540 544.320 ;
  LAYER metal2 ;
  RECT 1228.000 543.200 1231.540 544.320 ;
  LAYER metal1 ;
  RECT 1228.000 543.200 1231.540 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1160.420 543.200 1163.960 544.320 ;
  LAYER metal4 ;
  RECT 1160.420 543.200 1163.960 544.320 ;
  LAYER metal3 ;
  RECT 1160.420 543.200 1163.960 544.320 ;
  LAYER metal2 ;
  RECT 1160.420 543.200 1163.960 544.320 ;
  LAYER metal1 ;
  RECT 1160.420 543.200 1163.960 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1147.400 543.200 1150.940 544.320 ;
  LAYER metal4 ;
  RECT 1147.400 543.200 1150.940 544.320 ;
  LAYER metal3 ;
  RECT 1147.400 543.200 1150.940 544.320 ;
  LAYER metal2 ;
  RECT 1147.400 543.200 1150.940 544.320 ;
  LAYER metal1 ;
  RECT 1147.400 543.200 1150.940 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1133.760 543.200 1137.300 544.320 ;
  LAYER metal4 ;
  RECT 1133.760 543.200 1137.300 544.320 ;
  LAYER metal3 ;
  RECT 1133.760 543.200 1137.300 544.320 ;
  LAYER metal2 ;
  RECT 1133.760 543.200 1137.300 544.320 ;
  LAYER metal1 ;
  RECT 1133.760 543.200 1137.300 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1120.120 543.200 1123.660 544.320 ;
  LAYER metal4 ;
  RECT 1120.120 543.200 1123.660 544.320 ;
  LAYER metal3 ;
  RECT 1120.120 543.200 1123.660 544.320 ;
  LAYER metal2 ;
  RECT 1120.120 543.200 1123.660 544.320 ;
  LAYER metal1 ;
  RECT 1120.120 543.200 1123.660 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1107.100 543.200 1110.640 544.320 ;
  LAYER metal4 ;
  RECT 1107.100 543.200 1110.640 544.320 ;
  LAYER metal3 ;
  RECT 1107.100 543.200 1110.640 544.320 ;
  LAYER metal2 ;
  RECT 1107.100 543.200 1110.640 544.320 ;
  LAYER metal1 ;
  RECT 1107.100 543.200 1110.640 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1093.460 543.200 1097.000 544.320 ;
  LAYER metal4 ;
  RECT 1093.460 543.200 1097.000 544.320 ;
  LAYER metal3 ;
  RECT 1093.460 543.200 1097.000 544.320 ;
  LAYER metal2 ;
  RECT 1093.460 543.200 1097.000 544.320 ;
  LAYER metal1 ;
  RECT 1093.460 543.200 1097.000 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1025.880 543.200 1029.420 544.320 ;
  LAYER metal4 ;
  RECT 1025.880 543.200 1029.420 544.320 ;
  LAYER metal3 ;
  RECT 1025.880 543.200 1029.420 544.320 ;
  LAYER metal2 ;
  RECT 1025.880 543.200 1029.420 544.320 ;
  LAYER metal1 ;
  RECT 1025.880 543.200 1029.420 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1014.720 543.200 1018.260 544.320 ;
  LAYER metal4 ;
  RECT 1014.720 543.200 1018.260 544.320 ;
  LAYER metal3 ;
  RECT 1014.720 543.200 1018.260 544.320 ;
  LAYER metal2 ;
  RECT 1014.720 543.200 1018.260 544.320 ;
  LAYER metal1 ;
  RECT 1014.720 543.200 1018.260 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 999.220 543.200 1002.760 544.320 ;
  LAYER metal4 ;
  RECT 999.220 543.200 1002.760 544.320 ;
  LAYER metal3 ;
  RECT 999.220 543.200 1002.760 544.320 ;
  LAYER metal2 ;
  RECT 999.220 543.200 1002.760 544.320 ;
  LAYER metal1 ;
  RECT 999.220 543.200 1002.760 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 985.580 543.200 989.120 544.320 ;
  LAYER metal4 ;
  RECT 985.580 543.200 989.120 544.320 ;
  LAYER metal3 ;
  RECT 985.580 543.200 989.120 544.320 ;
  LAYER metal2 ;
  RECT 985.580 543.200 989.120 544.320 ;
  LAYER metal1 ;
  RECT 985.580 543.200 989.120 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 972.560 543.200 976.100 544.320 ;
  LAYER metal4 ;
  RECT 972.560 543.200 976.100 544.320 ;
  LAYER metal3 ;
  RECT 972.560 543.200 976.100 544.320 ;
  LAYER metal2 ;
  RECT 972.560 543.200 976.100 544.320 ;
  LAYER metal1 ;
  RECT 972.560 543.200 976.100 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 958.920 543.200 962.460 544.320 ;
  LAYER metal4 ;
  RECT 958.920 543.200 962.460 544.320 ;
  LAYER metal3 ;
  RECT 958.920 543.200 962.460 544.320 ;
  LAYER metal2 ;
  RECT 958.920 543.200 962.460 544.320 ;
  LAYER metal1 ;
  RECT 958.920 543.200 962.460 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 891.960 543.200 895.500 544.320 ;
  LAYER metal4 ;
  RECT 891.960 543.200 895.500 544.320 ;
  LAYER metal3 ;
  RECT 891.960 543.200 895.500 544.320 ;
  LAYER metal2 ;
  RECT 891.960 543.200 895.500 544.320 ;
  LAYER metal1 ;
  RECT 891.960 543.200 895.500 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 878.320 543.200 881.860 544.320 ;
  LAYER metal4 ;
  RECT 878.320 543.200 881.860 544.320 ;
  LAYER metal3 ;
  RECT 878.320 543.200 881.860 544.320 ;
  LAYER metal2 ;
  RECT 878.320 543.200 881.860 544.320 ;
  LAYER metal1 ;
  RECT 878.320 543.200 881.860 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 864.680 543.200 868.220 544.320 ;
  LAYER metal4 ;
  RECT 864.680 543.200 868.220 544.320 ;
  LAYER metal3 ;
  RECT 864.680 543.200 868.220 544.320 ;
  LAYER metal2 ;
  RECT 864.680 543.200 868.220 544.320 ;
  LAYER metal1 ;
  RECT 864.680 543.200 868.220 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 851.660 543.200 855.200 544.320 ;
  LAYER metal4 ;
  RECT 851.660 543.200 855.200 544.320 ;
  LAYER metal3 ;
  RECT 851.660 543.200 855.200 544.320 ;
  LAYER metal2 ;
  RECT 851.660 543.200 855.200 544.320 ;
  LAYER metal1 ;
  RECT 851.660 543.200 855.200 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 838.020 543.200 841.560 544.320 ;
  LAYER metal4 ;
  RECT 838.020 543.200 841.560 544.320 ;
  LAYER metal3 ;
  RECT 838.020 543.200 841.560 544.320 ;
  LAYER metal2 ;
  RECT 838.020 543.200 841.560 544.320 ;
  LAYER metal1 ;
  RECT 838.020 543.200 841.560 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 824.380 543.200 827.920 544.320 ;
  LAYER metal4 ;
  RECT 824.380 543.200 827.920 544.320 ;
  LAYER metal3 ;
  RECT 824.380 543.200 827.920 544.320 ;
  LAYER metal2 ;
  RECT 824.380 543.200 827.920 544.320 ;
  LAYER metal1 ;
  RECT 824.380 543.200 827.920 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 757.420 543.200 760.960 544.320 ;
  LAYER metal4 ;
  RECT 757.420 543.200 760.960 544.320 ;
  LAYER metal3 ;
  RECT 757.420 543.200 760.960 544.320 ;
  LAYER metal2 ;
  RECT 757.420 543.200 760.960 544.320 ;
  LAYER metal1 ;
  RECT 757.420 543.200 760.960 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 743.780 543.200 747.320 544.320 ;
  LAYER metal4 ;
  RECT 743.780 543.200 747.320 544.320 ;
  LAYER metal3 ;
  RECT 743.780 543.200 747.320 544.320 ;
  LAYER metal2 ;
  RECT 743.780 543.200 747.320 544.320 ;
  LAYER metal1 ;
  RECT 743.780 543.200 747.320 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 730.760 543.200 734.300 544.320 ;
  LAYER metal4 ;
  RECT 730.760 543.200 734.300 544.320 ;
  LAYER metal3 ;
  RECT 730.760 543.200 734.300 544.320 ;
  LAYER metal2 ;
  RECT 730.760 543.200 734.300 544.320 ;
  LAYER metal1 ;
  RECT 730.760 543.200 734.300 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 717.120 543.200 720.660 544.320 ;
  LAYER metal4 ;
  RECT 717.120 543.200 720.660 544.320 ;
  LAYER metal3 ;
  RECT 717.120 543.200 720.660 544.320 ;
  LAYER metal2 ;
  RECT 717.120 543.200 720.660 544.320 ;
  LAYER metal1 ;
  RECT 717.120 543.200 720.660 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 703.480 543.200 707.020 544.320 ;
  LAYER metal4 ;
  RECT 703.480 543.200 707.020 544.320 ;
  LAYER metal3 ;
  RECT 703.480 543.200 707.020 544.320 ;
  LAYER metal2 ;
  RECT 703.480 543.200 707.020 544.320 ;
  LAYER metal1 ;
  RECT 703.480 543.200 707.020 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 690.460 543.200 694.000 544.320 ;
  LAYER metal4 ;
  RECT 690.460 543.200 694.000 544.320 ;
  LAYER metal3 ;
  RECT 690.460 543.200 694.000 544.320 ;
  LAYER metal2 ;
  RECT 690.460 543.200 694.000 544.320 ;
  LAYER metal1 ;
  RECT 690.460 543.200 694.000 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 622.880 543.200 626.420 544.320 ;
  LAYER metal4 ;
  RECT 622.880 543.200 626.420 544.320 ;
  LAYER metal3 ;
  RECT 622.880 543.200 626.420 544.320 ;
  LAYER metal2 ;
  RECT 622.880 543.200 626.420 544.320 ;
  LAYER metal1 ;
  RECT 622.880 543.200 626.420 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 609.240 543.200 612.780 544.320 ;
  LAYER metal4 ;
  RECT 609.240 543.200 612.780 544.320 ;
  LAYER metal3 ;
  RECT 609.240 543.200 612.780 544.320 ;
  LAYER metal2 ;
  RECT 609.240 543.200 612.780 544.320 ;
  LAYER metal1 ;
  RECT 609.240 543.200 612.780 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 596.220 543.200 599.760 544.320 ;
  LAYER metal4 ;
  RECT 596.220 543.200 599.760 544.320 ;
  LAYER metal3 ;
  RECT 596.220 543.200 599.760 544.320 ;
  LAYER metal2 ;
  RECT 596.220 543.200 599.760 544.320 ;
  LAYER metal1 ;
  RECT 596.220 543.200 599.760 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 585.060 543.200 588.600 544.320 ;
  LAYER metal4 ;
  RECT 585.060 543.200 588.600 544.320 ;
  LAYER metal3 ;
  RECT 585.060 543.200 588.600 544.320 ;
  LAYER metal2 ;
  RECT 585.060 543.200 588.600 544.320 ;
  LAYER metal1 ;
  RECT 585.060 543.200 588.600 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 568.940 543.200 572.480 544.320 ;
  LAYER metal4 ;
  RECT 568.940 543.200 572.480 544.320 ;
  LAYER metal3 ;
  RECT 568.940 543.200 572.480 544.320 ;
  LAYER metal2 ;
  RECT 568.940 543.200 572.480 544.320 ;
  LAYER metal1 ;
  RECT 568.940 543.200 572.480 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 560.260 543.200 563.800 544.320 ;
  LAYER metal4 ;
  RECT 560.260 543.200 563.800 544.320 ;
  LAYER metal3 ;
  RECT 560.260 543.200 563.800 544.320 ;
  LAYER metal2 ;
  RECT 560.260 543.200 563.800 544.320 ;
  LAYER metal1 ;
  RECT 560.260 543.200 563.800 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 466.640 543.200 470.180 544.320 ;
  LAYER metal4 ;
  RECT 466.640 543.200 470.180 544.320 ;
  LAYER metal3 ;
  RECT 466.640 543.200 470.180 544.320 ;
  LAYER metal2 ;
  RECT 466.640 543.200 470.180 544.320 ;
  LAYER metal1 ;
  RECT 466.640 543.200 470.180 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 457.960 543.200 461.500 544.320 ;
  LAYER metal4 ;
  RECT 457.960 543.200 461.500 544.320 ;
  LAYER metal3 ;
  RECT 457.960 543.200 461.500 544.320 ;
  LAYER metal2 ;
  RECT 457.960 543.200 461.500 544.320 ;
  LAYER metal1 ;
  RECT 457.960 543.200 461.500 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 444.320 543.200 447.860 544.320 ;
  LAYER metal4 ;
  RECT 444.320 543.200 447.860 544.320 ;
  LAYER metal3 ;
  RECT 444.320 543.200 447.860 544.320 ;
  LAYER metal2 ;
  RECT 444.320 543.200 447.860 544.320 ;
  LAYER metal1 ;
  RECT 444.320 543.200 447.860 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 435.640 543.200 439.180 544.320 ;
  LAYER metal4 ;
  RECT 435.640 543.200 439.180 544.320 ;
  LAYER metal3 ;
  RECT 435.640 543.200 439.180 544.320 ;
  LAYER metal2 ;
  RECT 435.640 543.200 439.180 544.320 ;
  LAYER metal1 ;
  RECT 435.640 543.200 439.180 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 422.620 543.200 426.160 544.320 ;
  LAYER metal4 ;
  RECT 422.620 543.200 426.160 544.320 ;
  LAYER metal3 ;
  RECT 422.620 543.200 426.160 544.320 ;
  LAYER metal2 ;
  RECT 422.620 543.200 426.160 544.320 ;
  LAYER metal1 ;
  RECT 422.620 543.200 426.160 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 408.980 543.200 412.520 544.320 ;
  LAYER metal4 ;
  RECT 408.980 543.200 412.520 544.320 ;
  LAYER metal3 ;
  RECT 408.980 543.200 412.520 544.320 ;
  LAYER metal2 ;
  RECT 408.980 543.200 412.520 544.320 ;
  LAYER metal1 ;
  RECT 408.980 543.200 412.520 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 342.020 543.200 345.560 544.320 ;
  LAYER metal4 ;
  RECT 342.020 543.200 345.560 544.320 ;
  LAYER metal3 ;
  RECT 342.020 543.200 345.560 544.320 ;
  LAYER metal2 ;
  RECT 342.020 543.200 345.560 544.320 ;
  LAYER metal1 ;
  RECT 342.020 543.200 345.560 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 328.380 543.200 331.920 544.320 ;
  LAYER metal4 ;
  RECT 328.380 543.200 331.920 544.320 ;
  LAYER metal3 ;
  RECT 328.380 543.200 331.920 544.320 ;
  LAYER metal2 ;
  RECT 328.380 543.200 331.920 544.320 ;
  LAYER metal1 ;
  RECT 328.380 543.200 331.920 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 314.740 543.200 318.280 544.320 ;
  LAYER metal4 ;
  RECT 314.740 543.200 318.280 544.320 ;
  LAYER metal3 ;
  RECT 314.740 543.200 318.280 544.320 ;
  LAYER metal2 ;
  RECT 314.740 543.200 318.280 544.320 ;
  LAYER metal1 ;
  RECT 314.740 543.200 318.280 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 301.720 543.200 305.260 544.320 ;
  LAYER metal4 ;
  RECT 301.720 543.200 305.260 544.320 ;
  LAYER metal3 ;
  RECT 301.720 543.200 305.260 544.320 ;
  LAYER metal2 ;
  RECT 301.720 543.200 305.260 544.320 ;
  LAYER metal1 ;
  RECT 301.720 543.200 305.260 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 288.080 543.200 291.620 544.320 ;
  LAYER metal4 ;
  RECT 288.080 543.200 291.620 544.320 ;
  LAYER metal3 ;
  RECT 288.080 543.200 291.620 544.320 ;
  LAYER metal2 ;
  RECT 288.080 543.200 291.620 544.320 ;
  LAYER metal1 ;
  RECT 288.080 543.200 291.620 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 274.440 543.200 277.980 544.320 ;
  LAYER metal4 ;
  RECT 274.440 543.200 277.980 544.320 ;
  LAYER metal3 ;
  RECT 274.440 543.200 277.980 544.320 ;
  LAYER metal2 ;
  RECT 274.440 543.200 277.980 544.320 ;
  LAYER metal1 ;
  RECT 274.440 543.200 277.980 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 207.480 543.200 211.020 544.320 ;
  LAYER metal4 ;
  RECT 207.480 543.200 211.020 544.320 ;
  LAYER metal3 ;
  RECT 207.480 543.200 211.020 544.320 ;
  LAYER metal2 ;
  RECT 207.480 543.200 211.020 544.320 ;
  LAYER metal1 ;
  RECT 207.480 543.200 211.020 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 193.840 543.200 197.380 544.320 ;
  LAYER metal4 ;
  RECT 193.840 543.200 197.380 544.320 ;
  LAYER metal3 ;
  RECT 193.840 543.200 197.380 544.320 ;
  LAYER metal2 ;
  RECT 193.840 543.200 197.380 544.320 ;
  LAYER metal1 ;
  RECT 193.840 543.200 197.380 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 180.820 543.200 184.360 544.320 ;
  LAYER metal4 ;
  RECT 180.820 543.200 184.360 544.320 ;
  LAYER metal3 ;
  RECT 180.820 543.200 184.360 544.320 ;
  LAYER metal2 ;
  RECT 180.820 543.200 184.360 544.320 ;
  LAYER metal1 ;
  RECT 180.820 543.200 184.360 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 167.180 543.200 170.720 544.320 ;
  LAYER metal4 ;
  RECT 167.180 543.200 170.720 544.320 ;
  LAYER metal3 ;
  RECT 167.180 543.200 170.720 544.320 ;
  LAYER metal2 ;
  RECT 167.180 543.200 170.720 544.320 ;
  LAYER metal1 ;
  RECT 167.180 543.200 170.720 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 153.540 543.200 157.080 544.320 ;
  LAYER metal4 ;
  RECT 153.540 543.200 157.080 544.320 ;
  LAYER metal3 ;
  RECT 153.540 543.200 157.080 544.320 ;
  LAYER metal2 ;
  RECT 153.540 543.200 157.080 544.320 ;
  LAYER metal1 ;
  RECT 153.540 543.200 157.080 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 140.520 543.200 144.060 544.320 ;
  LAYER metal4 ;
  RECT 140.520 543.200 144.060 544.320 ;
  LAYER metal3 ;
  RECT 140.520 543.200 144.060 544.320 ;
  LAYER metal2 ;
  RECT 140.520 543.200 144.060 544.320 ;
  LAYER metal1 ;
  RECT 140.520 543.200 144.060 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 72.940 543.200 76.480 544.320 ;
  LAYER metal4 ;
  RECT 72.940 543.200 76.480 544.320 ;
  LAYER metal3 ;
  RECT 72.940 543.200 76.480 544.320 ;
  LAYER metal2 ;
  RECT 72.940 543.200 76.480 544.320 ;
  LAYER metal1 ;
  RECT 72.940 543.200 76.480 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 59.300 543.200 62.840 544.320 ;
  LAYER metal4 ;
  RECT 59.300 543.200 62.840 544.320 ;
  LAYER metal3 ;
  RECT 59.300 543.200 62.840 544.320 ;
  LAYER metal2 ;
  RECT 59.300 543.200 62.840 544.320 ;
  LAYER metal1 ;
  RECT 59.300 543.200 62.840 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 46.280 543.200 49.820 544.320 ;
  LAYER metal4 ;
  RECT 46.280 543.200 49.820 544.320 ;
  LAYER metal3 ;
  RECT 46.280 543.200 49.820 544.320 ;
  LAYER metal2 ;
  RECT 46.280 543.200 49.820 544.320 ;
  LAYER metal1 ;
  RECT 46.280 543.200 49.820 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 32.640 543.200 36.180 544.320 ;
  LAYER metal4 ;
  RECT 32.640 543.200 36.180 544.320 ;
  LAYER metal3 ;
  RECT 32.640 543.200 36.180 544.320 ;
  LAYER metal2 ;
  RECT 32.640 543.200 36.180 544.320 ;
  LAYER metal1 ;
  RECT 32.640 543.200 36.180 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 21.480 543.200 25.020 544.320 ;
  LAYER metal4 ;
  RECT 21.480 543.200 25.020 544.320 ;
  LAYER metal3 ;
  RECT 21.480 543.200 25.020 544.320 ;
  LAYER metal2 ;
  RECT 21.480 543.200 25.020 544.320 ;
  LAYER metal1 ;
  RECT 21.480 543.200 25.020 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 7.220 543.200 10.760 544.320 ;
  LAYER metal4 ;
  RECT 7.220 543.200 10.760 544.320 ;
  LAYER metal3 ;
  RECT 7.220 543.200 10.760 544.320 ;
  LAYER metal2 ;
  RECT 7.220 543.200 10.760 544.320 ;
  LAYER metal1 ;
  RECT 7.220 543.200 10.760 544.320 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1429.500 0.000 1433.040 1.120 ;
  LAYER metal4 ;
  RECT 1429.500 0.000 1433.040 1.120 ;
  LAYER metal3 ;
  RECT 1429.500 0.000 1433.040 1.120 ;
  LAYER metal2 ;
  RECT 1429.500 0.000 1433.040 1.120 ;
  LAYER metal1 ;
  RECT 1429.500 0.000 1433.040 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1415.860 0.000 1419.400 1.120 ;
  LAYER metal4 ;
  RECT 1415.860 0.000 1419.400 1.120 ;
  LAYER metal3 ;
  RECT 1415.860 0.000 1419.400 1.120 ;
  LAYER metal2 ;
  RECT 1415.860 0.000 1419.400 1.120 ;
  LAYER metal1 ;
  RECT 1415.860 0.000 1419.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1402.220 0.000 1405.760 1.120 ;
  LAYER metal4 ;
  RECT 1402.220 0.000 1405.760 1.120 ;
  LAYER metal3 ;
  RECT 1402.220 0.000 1405.760 1.120 ;
  LAYER metal2 ;
  RECT 1402.220 0.000 1405.760 1.120 ;
  LAYER metal1 ;
  RECT 1402.220 0.000 1405.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1389.200 0.000 1392.740 1.120 ;
  LAYER metal4 ;
  RECT 1389.200 0.000 1392.740 1.120 ;
  LAYER metal3 ;
  RECT 1389.200 0.000 1392.740 1.120 ;
  LAYER metal2 ;
  RECT 1389.200 0.000 1392.740 1.120 ;
  LAYER metal1 ;
  RECT 1389.200 0.000 1392.740 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1375.560 0.000 1379.100 1.120 ;
  LAYER metal4 ;
  RECT 1375.560 0.000 1379.100 1.120 ;
  LAYER metal3 ;
  RECT 1375.560 0.000 1379.100 1.120 ;
  LAYER metal2 ;
  RECT 1375.560 0.000 1379.100 1.120 ;
  LAYER metal1 ;
  RECT 1375.560 0.000 1379.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1361.920 0.000 1365.460 1.120 ;
  LAYER metal4 ;
  RECT 1361.920 0.000 1365.460 1.120 ;
  LAYER metal3 ;
  RECT 1361.920 0.000 1365.460 1.120 ;
  LAYER metal2 ;
  RECT 1361.920 0.000 1365.460 1.120 ;
  LAYER metal1 ;
  RECT 1361.920 0.000 1365.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1294.960 0.000 1298.500 1.120 ;
  LAYER metal4 ;
  RECT 1294.960 0.000 1298.500 1.120 ;
  LAYER metal3 ;
  RECT 1294.960 0.000 1298.500 1.120 ;
  LAYER metal2 ;
  RECT 1294.960 0.000 1298.500 1.120 ;
  LAYER metal1 ;
  RECT 1294.960 0.000 1298.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1281.320 0.000 1284.860 1.120 ;
  LAYER metal4 ;
  RECT 1281.320 0.000 1284.860 1.120 ;
  LAYER metal3 ;
  RECT 1281.320 0.000 1284.860 1.120 ;
  LAYER metal2 ;
  RECT 1281.320 0.000 1284.860 1.120 ;
  LAYER metal1 ;
  RECT 1281.320 0.000 1284.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1268.300 0.000 1271.840 1.120 ;
  LAYER metal4 ;
  RECT 1268.300 0.000 1271.840 1.120 ;
  LAYER metal3 ;
  RECT 1268.300 0.000 1271.840 1.120 ;
  LAYER metal2 ;
  RECT 1268.300 0.000 1271.840 1.120 ;
  LAYER metal1 ;
  RECT 1268.300 0.000 1271.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1254.660 0.000 1258.200 1.120 ;
  LAYER metal4 ;
  RECT 1254.660 0.000 1258.200 1.120 ;
  LAYER metal3 ;
  RECT 1254.660 0.000 1258.200 1.120 ;
  LAYER metal2 ;
  RECT 1254.660 0.000 1258.200 1.120 ;
  LAYER metal1 ;
  RECT 1254.660 0.000 1258.200 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1241.020 0.000 1244.560 1.120 ;
  LAYER metal4 ;
  RECT 1241.020 0.000 1244.560 1.120 ;
  LAYER metal3 ;
  RECT 1241.020 0.000 1244.560 1.120 ;
  LAYER metal2 ;
  RECT 1241.020 0.000 1244.560 1.120 ;
  LAYER metal1 ;
  RECT 1241.020 0.000 1244.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1228.000 0.000 1231.540 1.120 ;
  LAYER metal4 ;
  RECT 1228.000 0.000 1231.540 1.120 ;
  LAYER metal3 ;
  RECT 1228.000 0.000 1231.540 1.120 ;
  LAYER metal2 ;
  RECT 1228.000 0.000 1231.540 1.120 ;
  LAYER metal1 ;
  RECT 1228.000 0.000 1231.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1160.420 0.000 1163.960 1.120 ;
  LAYER metal4 ;
  RECT 1160.420 0.000 1163.960 1.120 ;
  LAYER metal3 ;
  RECT 1160.420 0.000 1163.960 1.120 ;
  LAYER metal2 ;
  RECT 1160.420 0.000 1163.960 1.120 ;
  LAYER metal1 ;
  RECT 1160.420 0.000 1163.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1147.400 0.000 1150.940 1.120 ;
  LAYER metal4 ;
  RECT 1147.400 0.000 1150.940 1.120 ;
  LAYER metal3 ;
  RECT 1147.400 0.000 1150.940 1.120 ;
  LAYER metal2 ;
  RECT 1147.400 0.000 1150.940 1.120 ;
  LAYER metal1 ;
  RECT 1147.400 0.000 1150.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1133.760 0.000 1137.300 1.120 ;
  LAYER metal4 ;
  RECT 1133.760 0.000 1137.300 1.120 ;
  LAYER metal3 ;
  RECT 1133.760 0.000 1137.300 1.120 ;
  LAYER metal2 ;
  RECT 1133.760 0.000 1137.300 1.120 ;
  LAYER metal1 ;
  RECT 1133.760 0.000 1137.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1120.120 0.000 1123.660 1.120 ;
  LAYER metal4 ;
  RECT 1120.120 0.000 1123.660 1.120 ;
  LAYER metal3 ;
  RECT 1120.120 0.000 1123.660 1.120 ;
  LAYER metal2 ;
  RECT 1120.120 0.000 1123.660 1.120 ;
  LAYER metal1 ;
  RECT 1120.120 0.000 1123.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1107.100 0.000 1110.640 1.120 ;
  LAYER metal4 ;
  RECT 1107.100 0.000 1110.640 1.120 ;
  LAYER metal3 ;
  RECT 1107.100 0.000 1110.640 1.120 ;
  LAYER metal2 ;
  RECT 1107.100 0.000 1110.640 1.120 ;
  LAYER metal1 ;
  RECT 1107.100 0.000 1110.640 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1093.460 0.000 1097.000 1.120 ;
  LAYER metal4 ;
  RECT 1093.460 0.000 1097.000 1.120 ;
  LAYER metal3 ;
  RECT 1093.460 0.000 1097.000 1.120 ;
  LAYER metal2 ;
  RECT 1093.460 0.000 1097.000 1.120 ;
  LAYER metal1 ;
  RECT 1093.460 0.000 1097.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1025.880 0.000 1029.420 1.120 ;
  LAYER metal4 ;
  RECT 1025.880 0.000 1029.420 1.120 ;
  LAYER metal3 ;
  RECT 1025.880 0.000 1029.420 1.120 ;
  LAYER metal2 ;
  RECT 1025.880 0.000 1029.420 1.120 ;
  LAYER metal1 ;
  RECT 1025.880 0.000 1029.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1014.720 0.000 1018.260 1.120 ;
  LAYER metal4 ;
  RECT 1014.720 0.000 1018.260 1.120 ;
  LAYER metal3 ;
  RECT 1014.720 0.000 1018.260 1.120 ;
  LAYER metal2 ;
  RECT 1014.720 0.000 1018.260 1.120 ;
  LAYER metal1 ;
  RECT 1014.720 0.000 1018.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 999.220 0.000 1002.760 1.120 ;
  LAYER metal4 ;
  RECT 999.220 0.000 1002.760 1.120 ;
  LAYER metal3 ;
  RECT 999.220 0.000 1002.760 1.120 ;
  LAYER metal2 ;
  RECT 999.220 0.000 1002.760 1.120 ;
  LAYER metal1 ;
  RECT 999.220 0.000 1002.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 985.580 0.000 989.120 1.120 ;
  LAYER metal4 ;
  RECT 985.580 0.000 989.120 1.120 ;
  LAYER metal3 ;
  RECT 985.580 0.000 989.120 1.120 ;
  LAYER metal2 ;
  RECT 985.580 0.000 989.120 1.120 ;
  LAYER metal1 ;
  RECT 985.580 0.000 989.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 972.560 0.000 976.100 1.120 ;
  LAYER metal4 ;
  RECT 972.560 0.000 976.100 1.120 ;
  LAYER metal3 ;
  RECT 972.560 0.000 976.100 1.120 ;
  LAYER metal2 ;
  RECT 972.560 0.000 976.100 1.120 ;
  LAYER metal1 ;
  RECT 972.560 0.000 976.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 958.920 0.000 962.460 1.120 ;
  LAYER metal4 ;
  RECT 958.920 0.000 962.460 1.120 ;
  LAYER metal3 ;
  RECT 958.920 0.000 962.460 1.120 ;
  LAYER metal2 ;
  RECT 958.920 0.000 962.460 1.120 ;
  LAYER metal1 ;
  RECT 958.920 0.000 962.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 891.960 0.000 895.500 1.120 ;
  LAYER metal4 ;
  RECT 891.960 0.000 895.500 1.120 ;
  LAYER metal3 ;
  RECT 891.960 0.000 895.500 1.120 ;
  LAYER metal2 ;
  RECT 891.960 0.000 895.500 1.120 ;
  LAYER metal1 ;
  RECT 891.960 0.000 895.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 878.320 0.000 881.860 1.120 ;
  LAYER metal4 ;
  RECT 878.320 0.000 881.860 1.120 ;
  LAYER metal3 ;
  RECT 878.320 0.000 881.860 1.120 ;
  LAYER metal2 ;
  RECT 878.320 0.000 881.860 1.120 ;
  LAYER metal1 ;
  RECT 878.320 0.000 881.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 864.680 0.000 868.220 1.120 ;
  LAYER metal4 ;
  RECT 864.680 0.000 868.220 1.120 ;
  LAYER metal3 ;
  RECT 864.680 0.000 868.220 1.120 ;
  LAYER metal2 ;
  RECT 864.680 0.000 868.220 1.120 ;
  LAYER metal1 ;
  RECT 864.680 0.000 868.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 851.660 0.000 855.200 1.120 ;
  LAYER metal4 ;
  RECT 851.660 0.000 855.200 1.120 ;
  LAYER metal3 ;
  RECT 851.660 0.000 855.200 1.120 ;
  LAYER metal2 ;
  RECT 851.660 0.000 855.200 1.120 ;
  LAYER metal1 ;
  RECT 851.660 0.000 855.200 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 838.020 0.000 841.560 1.120 ;
  LAYER metal4 ;
  RECT 838.020 0.000 841.560 1.120 ;
  LAYER metal3 ;
  RECT 838.020 0.000 841.560 1.120 ;
  LAYER metal2 ;
  RECT 838.020 0.000 841.560 1.120 ;
  LAYER metal1 ;
  RECT 838.020 0.000 841.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 824.380 0.000 827.920 1.120 ;
  LAYER metal4 ;
  RECT 824.380 0.000 827.920 1.120 ;
  LAYER metal3 ;
  RECT 824.380 0.000 827.920 1.120 ;
  LAYER metal2 ;
  RECT 824.380 0.000 827.920 1.120 ;
  LAYER metal1 ;
  RECT 824.380 0.000 827.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 757.420 0.000 760.960 1.120 ;
  LAYER metal4 ;
  RECT 757.420 0.000 760.960 1.120 ;
  LAYER metal3 ;
  RECT 757.420 0.000 760.960 1.120 ;
  LAYER metal2 ;
  RECT 757.420 0.000 760.960 1.120 ;
  LAYER metal1 ;
  RECT 757.420 0.000 760.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 743.780 0.000 747.320 1.120 ;
  LAYER metal4 ;
  RECT 743.780 0.000 747.320 1.120 ;
  LAYER metal3 ;
  RECT 743.780 0.000 747.320 1.120 ;
  LAYER metal2 ;
  RECT 743.780 0.000 747.320 1.120 ;
  LAYER metal1 ;
  RECT 743.780 0.000 747.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 730.760 0.000 734.300 1.120 ;
  LAYER metal4 ;
  RECT 730.760 0.000 734.300 1.120 ;
  LAYER metal3 ;
  RECT 730.760 0.000 734.300 1.120 ;
  LAYER metal2 ;
  RECT 730.760 0.000 734.300 1.120 ;
  LAYER metal1 ;
  RECT 730.760 0.000 734.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 717.120 0.000 720.660 1.120 ;
  LAYER metal4 ;
  RECT 717.120 0.000 720.660 1.120 ;
  LAYER metal3 ;
  RECT 717.120 0.000 720.660 1.120 ;
  LAYER metal2 ;
  RECT 717.120 0.000 720.660 1.120 ;
  LAYER metal1 ;
  RECT 717.120 0.000 720.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 703.480 0.000 707.020 1.120 ;
  LAYER metal4 ;
  RECT 703.480 0.000 707.020 1.120 ;
  LAYER metal3 ;
  RECT 703.480 0.000 707.020 1.120 ;
  LAYER metal2 ;
  RECT 703.480 0.000 707.020 1.120 ;
  LAYER metal1 ;
  RECT 703.480 0.000 707.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 690.460 0.000 694.000 1.120 ;
  LAYER metal4 ;
  RECT 690.460 0.000 694.000 1.120 ;
  LAYER metal3 ;
  RECT 690.460 0.000 694.000 1.120 ;
  LAYER metal2 ;
  RECT 690.460 0.000 694.000 1.120 ;
  LAYER metal1 ;
  RECT 690.460 0.000 694.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 622.880 0.000 626.420 1.120 ;
  LAYER metal4 ;
  RECT 622.880 0.000 626.420 1.120 ;
  LAYER metal3 ;
  RECT 622.880 0.000 626.420 1.120 ;
  LAYER metal2 ;
  RECT 622.880 0.000 626.420 1.120 ;
  LAYER metal1 ;
  RECT 622.880 0.000 626.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 609.240 0.000 612.780 1.120 ;
  LAYER metal4 ;
  RECT 609.240 0.000 612.780 1.120 ;
  LAYER metal3 ;
  RECT 609.240 0.000 612.780 1.120 ;
  LAYER metal2 ;
  RECT 609.240 0.000 612.780 1.120 ;
  LAYER metal1 ;
  RECT 609.240 0.000 612.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 596.220 0.000 599.760 1.120 ;
  LAYER metal4 ;
  RECT 596.220 0.000 599.760 1.120 ;
  LAYER metal3 ;
  RECT 596.220 0.000 599.760 1.120 ;
  LAYER metal2 ;
  RECT 596.220 0.000 599.760 1.120 ;
  LAYER metal1 ;
  RECT 596.220 0.000 599.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 585.060 0.000 588.600 1.120 ;
  LAYER metal4 ;
  RECT 585.060 0.000 588.600 1.120 ;
  LAYER metal3 ;
  RECT 585.060 0.000 588.600 1.120 ;
  LAYER metal2 ;
  RECT 585.060 0.000 588.600 1.120 ;
  LAYER metal1 ;
  RECT 585.060 0.000 588.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 568.940 0.000 572.480 1.120 ;
  LAYER metal4 ;
  RECT 568.940 0.000 572.480 1.120 ;
  LAYER metal3 ;
  RECT 568.940 0.000 572.480 1.120 ;
  LAYER metal2 ;
  RECT 568.940 0.000 572.480 1.120 ;
  LAYER metal1 ;
  RECT 568.940 0.000 572.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 560.260 0.000 563.800 1.120 ;
  LAYER metal4 ;
  RECT 560.260 0.000 563.800 1.120 ;
  LAYER metal3 ;
  RECT 560.260 0.000 563.800 1.120 ;
  LAYER metal2 ;
  RECT 560.260 0.000 563.800 1.120 ;
  LAYER metal1 ;
  RECT 560.260 0.000 563.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 466.640 0.000 470.180 1.120 ;
  LAYER metal4 ;
  RECT 466.640 0.000 470.180 1.120 ;
  LAYER metal3 ;
  RECT 466.640 0.000 470.180 1.120 ;
  LAYER metal2 ;
  RECT 466.640 0.000 470.180 1.120 ;
  LAYER metal1 ;
  RECT 466.640 0.000 470.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 457.960 0.000 461.500 1.120 ;
  LAYER metal4 ;
  RECT 457.960 0.000 461.500 1.120 ;
  LAYER metal3 ;
  RECT 457.960 0.000 461.500 1.120 ;
  LAYER metal2 ;
  RECT 457.960 0.000 461.500 1.120 ;
  LAYER metal1 ;
  RECT 457.960 0.000 461.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 444.320 0.000 447.860 1.120 ;
  LAYER metal4 ;
  RECT 444.320 0.000 447.860 1.120 ;
  LAYER metal3 ;
  RECT 444.320 0.000 447.860 1.120 ;
  LAYER metal2 ;
  RECT 444.320 0.000 447.860 1.120 ;
  LAYER metal1 ;
  RECT 444.320 0.000 447.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER metal4 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER metal3 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER metal2 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER metal1 ;
  RECT 435.640 0.000 439.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 422.620 0.000 426.160 1.120 ;
  LAYER metal4 ;
  RECT 422.620 0.000 426.160 1.120 ;
  LAYER metal3 ;
  RECT 422.620 0.000 426.160 1.120 ;
  LAYER metal2 ;
  RECT 422.620 0.000 426.160 1.120 ;
  LAYER metal1 ;
  RECT 422.620 0.000 426.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 408.980 0.000 412.520 1.120 ;
  LAYER metal4 ;
  RECT 408.980 0.000 412.520 1.120 ;
  LAYER metal3 ;
  RECT 408.980 0.000 412.520 1.120 ;
  LAYER metal2 ;
  RECT 408.980 0.000 412.520 1.120 ;
  LAYER metal1 ;
  RECT 408.980 0.000 412.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 342.020 0.000 345.560 1.120 ;
  LAYER metal4 ;
  RECT 342.020 0.000 345.560 1.120 ;
  LAYER metal3 ;
  RECT 342.020 0.000 345.560 1.120 ;
  LAYER metal2 ;
  RECT 342.020 0.000 345.560 1.120 ;
  LAYER metal1 ;
  RECT 342.020 0.000 345.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER metal4 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER metal3 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER metal2 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER metal1 ;
  RECT 328.380 0.000 331.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 314.740 0.000 318.280 1.120 ;
  LAYER metal4 ;
  RECT 314.740 0.000 318.280 1.120 ;
  LAYER metal3 ;
  RECT 314.740 0.000 318.280 1.120 ;
  LAYER metal2 ;
  RECT 314.740 0.000 318.280 1.120 ;
  LAYER metal1 ;
  RECT 314.740 0.000 318.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 301.720 0.000 305.260 1.120 ;
  LAYER metal4 ;
  RECT 301.720 0.000 305.260 1.120 ;
  LAYER metal3 ;
  RECT 301.720 0.000 305.260 1.120 ;
  LAYER metal2 ;
  RECT 301.720 0.000 305.260 1.120 ;
  LAYER metal1 ;
  RECT 301.720 0.000 305.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 288.080 0.000 291.620 1.120 ;
  LAYER metal4 ;
  RECT 288.080 0.000 291.620 1.120 ;
  LAYER metal3 ;
  RECT 288.080 0.000 291.620 1.120 ;
  LAYER metal2 ;
  RECT 288.080 0.000 291.620 1.120 ;
  LAYER metal1 ;
  RECT 288.080 0.000 291.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER metal4 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER metal3 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER metal2 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER metal1 ;
  RECT 274.440 0.000 277.980 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 207.480 0.000 211.020 1.120 ;
  LAYER metal4 ;
  RECT 207.480 0.000 211.020 1.120 ;
  LAYER metal3 ;
  RECT 207.480 0.000 211.020 1.120 ;
  LAYER metal2 ;
  RECT 207.480 0.000 211.020 1.120 ;
  LAYER metal1 ;
  RECT 207.480 0.000 211.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 193.840 0.000 197.380 1.120 ;
  LAYER metal4 ;
  RECT 193.840 0.000 197.380 1.120 ;
  LAYER metal3 ;
  RECT 193.840 0.000 197.380 1.120 ;
  LAYER metal2 ;
  RECT 193.840 0.000 197.380 1.120 ;
  LAYER metal1 ;
  RECT 193.840 0.000 197.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 180.820 0.000 184.360 1.120 ;
  LAYER metal4 ;
  RECT 180.820 0.000 184.360 1.120 ;
  LAYER metal3 ;
  RECT 180.820 0.000 184.360 1.120 ;
  LAYER metal2 ;
  RECT 180.820 0.000 184.360 1.120 ;
  LAYER metal1 ;
  RECT 180.820 0.000 184.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 167.180 0.000 170.720 1.120 ;
  LAYER metal4 ;
  RECT 167.180 0.000 170.720 1.120 ;
  LAYER metal3 ;
  RECT 167.180 0.000 170.720 1.120 ;
  LAYER metal2 ;
  RECT 167.180 0.000 170.720 1.120 ;
  LAYER metal1 ;
  RECT 167.180 0.000 170.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 153.540 0.000 157.080 1.120 ;
  LAYER metal4 ;
  RECT 153.540 0.000 157.080 1.120 ;
  LAYER metal3 ;
  RECT 153.540 0.000 157.080 1.120 ;
  LAYER metal2 ;
  RECT 153.540 0.000 157.080 1.120 ;
  LAYER metal1 ;
  RECT 153.540 0.000 157.080 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER metal4 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER metal3 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER metal2 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER metal1 ;
  RECT 140.520 0.000 144.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 72.940 0.000 76.480 1.120 ;
  LAYER metal4 ;
  RECT 72.940 0.000 76.480 1.120 ;
  LAYER metal3 ;
  RECT 72.940 0.000 76.480 1.120 ;
  LAYER metal2 ;
  RECT 72.940 0.000 76.480 1.120 ;
  LAYER metal1 ;
  RECT 72.940 0.000 76.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER metal4 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER metal3 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER metal2 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER metal1 ;
  RECT 59.300 0.000 62.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER metal4 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER metal3 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER metal2 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER metal1 ;
  RECT 46.280 0.000 49.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER metal4 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER metal3 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER metal2 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER metal1 ;
  RECT 32.640 0.000 36.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 21.480 0.000 25.020 1.120 ;
  LAYER metal4 ;
  RECT 21.480 0.000 25.020 1.120 ;
  LAYER metal3 ;
  RECT 21.480 0.000 25.020 1.120 ;
  LAYER metal2 ;
  RECT 21.480 0.000 25.020 1.120 ;
  LAYER metal1 ;
  RECT 21.480 0.000 25.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER metal4 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER metal3 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER metal2 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER metal1 ;
  RECT 7.220 0.000 10.760 1.120 ;
 END
END VCC
PIN DIB47
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1422.960 543.200 1424.080 544.320 ;
  LAYER metal4 ;
  RECT 1422.960 543.200 1424.080 544.320 ;
  LAYER metal3 ;
  RECT 1422.960 543.200 1424.080 544.320 ;
  LAYER metal2 ;
  RECT 1422.960 543.200 1424.080 544.320 ;
  LAYER metal1 ;
  RECT 1422.960 543.200 1424.080 544.320 ;
 END
END DIB47
PIN DOB47
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1409.320 543.200 1410.440 544.320 ;
  LAYER metal4 ;
  RECT 1409.320 543.200 1410.440 544.320 ;
  LAYER metal3 ;
  RECT 1409.320 543.200 1410.440 544.320 ;
  LAYER metal2 ;
  RECT 1409.320 543.200 1410.440 544.320 ;
  LAYER metal1 ;
  RECT 1409.320 543.200 1410.440 544.320 ;
 END
END DOB47
PIN DIB46
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1395.680 543.200 1396.800 544.320 ;
  LAYER metal4 ;
  RECT 1395.680 543.200 1396.800 544.320 ;
  LAYER metal3 ;
  RECT 1395.680 543.200 1396.800 544.320 ;
  LAYER metal2 ;
  RECT 1395.680 543.200 1396.800 544.320 ;
  LAYER metal1 ;
  RECT 1395.680 543.200 1396.800 544.320 ;
 END
END DIB46
PIN DOB46
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1382.660 543.200 1383.780 544.320 ;
  LAYER metal4 ;
  RECT 1382.660 543.200 1383.780 544.320 ;
  LAYER metal3 ;
  RECT 1382.660 543.200 1383.780 544.320 ;
  LAYER metal2 ;
  RECT 1382.660 543.200 1383.780 544.320 ;
  LAYER metal1 ;
  RECT 1382.660 543.200 1383.780 544.320 ;
 END
END DOB46
PIN DIB45
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1369.020 543.200 1370.140 544.320 ;
  LAYER metal4 ;
  RECT 1369.020 543.200 1370.140 544.320 ;
  LAYER metal3 ;
  RECT 1369.020 543.200 1370.140 544.320 ;
  LAYER metal2 ;
  RECT 1369.020 543.200 1370.140 544.320 ;
  LAYER metal1 ;
  RECT 1369.020 543.200 1370.140 544.320 ;
 END
END DIB45
PIN DOB45
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1355.380 543.200 1356.500 544.320 ;
  LAYER metal4 ;
  RECT 1355.380 543.200 1356.500 544.320 ;
  LAYER metal3 ;
  RECT 1355.380 543.200 1356.500 544.320 ;
  LAYER metal2 ;
  RECT 1355.380 543.200 1356.500 544.320 ;
  LAYER metal1 ;
  RECT 1355.380 543.200 1356.500 544.320 ;
 END
END DOB45
PIN DIB44
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1342.360 543.200 1343.480 544.320 ;
  LAYER metal4 ;
  RECT 1342.360 543.200 1343.480 544.320 ;
  LAYER metal3 ;
  RECT 1342.360 543.200 1343.480 544.320 ;
  LAYER metal2 ;
  RECT 1342.360 543.200 1343.480 544.320 ;
  LAYER metal1 ;
  RECT 1342.360 543.200 1343.480 544.320 ;
 END
END DIB44
PIN DOB44
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1328.720 543.200 1329.840 544.320 ;
  LAYER metal4 ;
  RECT 1328.720 543.200 1329.840 544.320 ;
  LAYER metal3 ;
  RECT 1328.720 543.200 1329.840 544.320 ;
  LAYER metal2 ;
  RECT 1328.720 543.200 1329.840 544.320 ;
  LAYER metal1 ;
  RECT 1328.720 543.200 1329.840 544.320 ;
 END
END DOB44
PIN DIB43
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1315.080 543.200 1316.200 544.320 ;
  LAYER metal4 ;
  RECT 1315.080 543.200 1316.200 544.320 ;
  LAYER metal3 ;
  RECT 1315.080 543.200 1316.200 544.320 ;
  LAYER metal2 ;
  RECT 1315.080 543.200 1316.200 544.320 ;
  LAYER metal1 ;
  RECT 1315.080 543.200 1316.200 544.320 ;
 END
END DIB43
PIN DOB43
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1302.060 543.200 1303.180 544.320 ;
  LAYER metal4 ;
  RECT 1302.060 543.200 1303.180 544.320 ;
  LAYER metal3 ;
  RECT 1302.060 543.200 1303.180 544.320 ;
  LAYER metal2 ;
  RECT 1302.060 543.200 1303.180 544.320 ;
  LAYER metal1 ;
  RECT 1302.060 543.200 1303.180 544.320 ;
 END
END DOB43
PIN DIB42
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1288.420 543.200 1289.540 544.320 ;
  LAYER metal4 ;
  RECT 1288.420 543.200 1289.540 544.320 ;
  LAYER metal3 ;
  RECT 1288.420 543.200 1289.540 544.320 ;
  LAYER metal2 ;
  RECT 1288.420 543.200 1289.540 544.320 ;
  LAYER metal1 ;
  RECT 1288.420 543.200 1289.540 544.320 ;
 END
END DIB42
PIN DOB42
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1274.780 543.200 1275.900 544.320 ;
  LAYER metal4 ;
  RECT 1274.780 543.200 1275.900 544.320 ;
  LAYER metal3 ;
  RECT 1274.780 543.200 1275.900 544.320 ;
  LAYER metal2 ;
  RECT 1274.780 543.200 1275.900 544.320 ;
  LAYER metal1 ;
  RECT 1274.780 543.200 1275.900 544.320 ;
 END
END DOB42
PIN DIB41
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1261.760 543.200 1262.880 544.320 ;
  LAYER metal4 ;
  RECT 1261.760 543.200 1262.880 544.320 ;
  LAYER metal3 ;
  RECT 1261.760 543.200 1262.880 544.320 ;
  LAYER metal2 ;
  RECT 1261.760 543.200 1262.880 544.320 ;
  LAYER metal1 ;
  RECT 1261.760 543.200 1262.880 544.320 ;
 END
END DIB41
PIN DOB41
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1248.120 543.200 1249.240 544.320 ;
  LAYER metal4 ;
  RECT 1248.120 543.200 1249.240 544.320 ;
  LAYER metal3 ;
  RECT 1248.120 543.200 1249.240 544.320 ;
  LAYER metal2 ;
  RECT 1248.120 543.200 1249.240 544.320 ;
  LAYER metal1 ;
  RECT 1248.120 543.200 1249.240 544.320 ;
 END
END DOB41
PIN DIB40
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1234.480 543.200 1235.600 544.320 ;
  LAYER metal4 ;
  RECT 1234.480 543.200 1235.600 544.320 ;
  LAYER metal3 ;
  RECT 1234.480 543.200 1235.600 544.320 ;
  LAYER metal2 ;
  RECT 1234.480 543.200 1235.600 544.320 ;
  LAYER metal1 ;
  RECT 1234.480 543.200 1235.600 544.320 ;
 END
END DIB40
PIN DOB40
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1221.460 543.200 1222.580 544.320 ;
  LAYER metal4 ;
  RECT 1221.460 543.200 1222.580 544.320 ;
  LAYER metal3 ;
  RECT 1221.460 543.200 1222.580 544.320 ;
  LAYER metal2 ;
  RECT 1221.460 543.200 1222.580 544.320 ;
  LAYER metal1 ;
  RECT 1221.460 543.200 1222.580 544.320 ;
 END
END DOB40
PIN DIB39
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1207.820 543.200 1208.940 544.320 ;
  LAYER metal4 ;
  RECT 1207.820 543.200 1208.940 544.320 ;
  LAYER metal3 ;
  RECT 1207.820 543.200 1208.940 544.320 ;
  LAYER metal2 ;
  RECT 1207.820 543.200 1208.940 544.320 ;
  LAYER metal1 ;
  RECT 1207.820 543.200 1208.940 544.320 ;
 END
END DIB39
PIN DOB39
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1194.180 543.200 1195.300 544.320 ;
  LAYER metal4 ;
  RECT 1194.180 543.200 1195.300 544.320 ;
  LAYER metal3 ;
  RECT 1194.180 543.200 1195.300 544.320 ;
  LAYER metal2 ;
  RECT 1194.180 543.200 1195.300 544.320 ;
  LAYER metal1 ;
  RECT 1194.180 543.200 1195.300 544.320 ;
 END
END DOB39
PIN DIB38
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1181.160 543.200 1182.280 544.320 ;
  LAYER metal4 ;
  RECT 1181.160 543.200 1182.280 544.320 ;
  LAYER metal3 ;
  RECT 1181.160 543.200 1182.280 544.320 ;
  LAYER metal2 ;
  RECT 1181.160 543.200 1182.280 544.320 ;
  LAYER metal1 ;
  RECT 1181.160 543.200 1182.280 544.320 ;
 END
END DIB38
PIN DOB38
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1167.520 543.200 1168.640 544.320 ;
  LAYER metal4 ;
  RECT 1167.520 543.200 1168.640 544.320 ;
  LAYER metal3 ;
  RECT 1167.520 543.200 1168.640 544.320 ;
  LAYER metal2 ;
  RECT 1167.520 543.200 1168.640 544.320 ;
  LAYER metal1 ;
  RECT 1167.520 543.200 1168.640 544.320 ;
 END
END DOB38
PIN DIB37
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1153.880 543.200 1155.000 544.320 ;
  LAYER metal4 ;
  RECT 1153.880 543.200 1155.000 544.320 ;
  LAYER metal3 ;
  RECT 1153.880 543.200 1155.000 544.320 ;
  LAYER metal2 ;
  RECT 1153.880 543.200 1155.000 544.320 ;
  LAYER metal1 ;
  RECT 1153.880 543.200 1155.000 544.320 ;
 END
END DIB37
PIN DOB37
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1140.860 543.200 1141.980 544.320 ;
  LAYER metal4 ;
  RECT 1140.860 543.200 1141.980 544.320 ;
  LAYER metal3 ;
  RECT 1140.860 543.200 1141.980 544.320 ;
  LAYER metal2 ;
  RECT 1140.860 543.200 1141.980 544.320 ;
  LAYER metal1 ;
  RECT 1140.860 543.200 1141.980 544.320 ;
 END
END DOB37
PIN DIB36
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1127.220 543.200 1128.340 544.320 ;
  LAYER metal4 ;
  RECT 1127.220 543.200 1128.340 544.320 ;
  LAYER metal3 ;
  RECT 1127.220 543.200 1128.340 544.320 ;
  LAYER metal2 ;
  RECT 1127.220 543.200 1128.340 544.320 ;
  LAYER metal1 ;
  RECT 1127.220 543.200 1128.340 544.320 ;
 END
END DIB36
PIN DOB36
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1113.580 543.200 1114.700 544.320 ;
  LAYER metal4 ;
  RECT 1113.580 543.200 1114.700 544.320 ;
  LAYER metal3 ;
  RECT 1113.580 543.200 1114.700 544.320 ;
  LAYER metal2 ;
  RECT 1113.580 543.200 1114.700 544.320 ;
  LAYER metal1 ;
  RECT 1113.580 543.200 1114.700 544.320 ;
 END
END DOB36
PIN DIB35
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1100.560 543.200 1101.680 544.320 ;
  LAYER metal4 ;
  RECT 1100.560 543.200 1101.680 544.320 ;
  LAYER metal3 ;
  RECT 1100.560 543.200 1101.680 544.320 ;
  LAYER metal2 ;
  RECT 1100.560 543.200 1101.680 544.320 ;
  LAYER metal1 ;
  RECT 1100.560 543.200 1101.680 544.320 ;
 END
END DIB35
PIN DOB35
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1086.920 543.200 1088.040 544.320 ;
  LAYER metal4 ;
  RECT 1086.920 543.200 1088.040 544.320 ;
  LAYER metal3 ;
  RECT 1086.920 543.200 1088.040 544.320 ;
  LAYER metal2 ;
  RECT 1086.920 543.200 1088.040 544.320 ;
  LAYER metal1 ;
  RECT 1086.920 543.200 1088.040 544.320 ;
 END
END DOB35
PIN DIB34
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1073.280 543.200 1074.400 544.320 ;
  LAYER metal4 ;
  RECT 1073.280 543.200 1074.400 544.320 ;
  LAYER metal3 ;
  RECT 1073.280 543.200 1074.400 544.320 ;
  LAYER metal2 ;
  RECT 1073.280 543.200 1074.400 544.320 ;
  LAYER metal1 ;
  RECT 1073.280 543.200 1074.400 544.320 ;
 END
END DIB34
PIN DOB34
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1059.640 543.200 1060.760 544.320 ;
  LAYER metal4 ;
  RECT 1059.640 543.200 1060.760 544.320 ;
  LAYER metal3 ;
  RECT 1059.640 543.200 1060.760 544.320 ;
  LAYER metal2 ;
  RECT 1059.640 543.200 1060.760 544.320 ;
  LAYER metal1 ;
  RECT 1059.640 543.200 1060.760 544.320 ;
 END
END DOB34
PIN DIB33
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1046.620 543.200 1047.740 544.320 ;
  LAYER metal4 ;
  RECT 1046.620 543.200 1047.740 544.320 ;
  LAYER metal3 ;
  RECT 1046.620 543.200 1047.740 544.320 ;
  LAYER metal2 ;
  RECT 1046.620 543.200 1047.740 544.320 ;
  LAYER metal1 ;
  RECT 1046.620 543.200 1047.740 544.320 ;
 END
END DIB33
PIN DOB33
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1032.980 543.200 1034.100 544.320 ;
  LAYER metal4 ;
  RECT 1032.980 543.200 1034.100 544.320 ;
  LAYER metal3 ;
  RECT 1032.980 543.200 1034.100 544.320 ;
  LAYER metal2 ;
  RECT 1032.980 543.200 1034.100 544.320 ;
  LAYER metal1 ;
  RECT 1032.980 543.200 1034.100 544.320 ;
 END
END DOB33
PIN DIB32
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1019.340 543.200 1020.460 544.320 ;
  LAYER metal4 ;
  RECT 1019.340 543.200 1020.460 544.320 ;
  LAYER metal3 ;
  RECT 1019.340 543.200 1020.460 544.320 ;
  LAYER metal2 ;
  RECT 1019.340 543.200 1020.460 544.320 ;
  LAYER metal1 ;
  RECT 1019.340 543.200 1020.460 544.320 ;
 END
END DIB32
PIN WEBN2
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1008.180 543.200 1009.300 544.320 ;
  LAYER metal4 ;
  RECT 1008.180 543.200 1009.300 544.320 ;
  LAYER metal3 ;
  RECT 1008.180 543.200 1009.300 544.320 ;
  LAYER metal2 ;
  RECT 1008.180 543.200 1009.300 544.320 ;
  LAYER metal1 ;
  RECT 1008.180 543.200 1009.300 544.320 ;
 END
END WEBN2
PIN DOB32
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1006.320 543.200 1007.440 544.320 ;
  LAYER metal4 ;
  RECT 1006.320 543.200 1007.440 544.320 ;
  LAYER metal3 ;
  RECT 1006.320 543.200 1007.440 544.320 ;
  LAYER metal2 ;
  RECT 1006.320 543.200 1007.440 544.320 ;
  LAYER metal1 ;
  RECT 1006.320 543.200 1007.440 544.320 ;
 END
END DOB32
PIN DIB31
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 992.680 543.200 993.800 544.320 ;
  LAYER metal4 ;
  RECT 992.680 543.200 993.800 544.320 ;
  LAYER metal3 ;
  RECT 992.680 543.200 993.800 544.320 ;
  LAYER metal2 ;
  RECT 992.680 543.200 993.800 544.320 ;
  LAYER metal1 ;
  RECT 992.680 543.200 993.800 544.320 ;
 END
END DIB31
PIN DOB31
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 979.040 543.200 980.160 544.320 ;
  LAYER metal4 ;
  RECT 979.040 543.200 980.160 544.320 ;
  LAYER metal3 ;
  RECT 979.040 543.200 980.160 544.320 ;
  LAYER metal2 ;
  RECT 979.040 543.200 980.160 544.320 ;
  LAYER metal1 ;
  RECT 979.040 543.200 980.160 544.320 ;
 END
END DOB31
PIN DIB30
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 966.020 543.200 967.140 544.320 ;
  LAYER metal4 ;
  RECT 966.020 543.200 967.140 544.320 ;
  LAYER metal3 ;
  RECT 966.020 543.200 967.140 544.320 ;
  LAYER metal2 ;
  RECT 966.020 543.200 967.140 544.320 ;
  LAYER metal1 ;
  RECT 966.020 543.200 967.140 544.320 ;
 END
END DIB30
PIN DOB30
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 952.380 543.200 953.500 544.320 ;
  LAYER metal4 ;
  RECT 952.380 543.200 953.500 544.320 ;
  LAYER metal3 ;
  RECT 952.380 543.200 953.500 544.320 ;
  LAYER metal2 ;
  RECT 952.380 543.200 953.500 544.320 ;
  LAYER metal1 ;
  RECT 952.380 543.200 953.500 544.320 ;
 END
END DOB30
PIN DIB29
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 938.740 543.200 939.860 544.320 ;
  LAYER metal4 ;
  RECT 938.740 543.200 939.860 544.320 ;
  LAYER metal3 ;
  RECT 938.740 543.200 939.860 544.320 ;
  LAYER metal2 ;
  RECT 938.740 543.200 939.860 544.320 ;
  LAYER metal1 ;
  RECT 938.740 543.200 939.860 544.320 ;
 END
END DIB29
PIN DOB29
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 925.720 543.200 926.840 544.320 ;
  LAYER metal4 ;
  RECT 925.720 543.200 926.840 544.320 ;
  LAYER metal3 ;
  RECT 925.720 543.200 926.840 544.320 ;
  LAYER metal2 ;
  RECT 925.720 543.200 926.840 544.320 ;
  LAYER metal1 ;
  RECT 925.720 543.200 926.840 544.320 ;
 END
END DOB29
PIN DIB28
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 912.080 543.200 913.200 544.320 ;
  LAYER metal4 ;
  RECT 912.080 543.200 913.200 544.320 ;
  LAYER metal3 ;
  RECT 912.080 543.200 913.200 544.320 ;
  LAYER metal2 ;
  RECT 912.080 543.200 913.200 544.320 ;
  LAYER metal1 ;
  RECT 912.080 543.200 913.200 544.320 ;
 END
END DIB28
PIN DOB28
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 898.440 543.200 899.560 544.320 ;
  LAYER metal4 ;
  RECT 898.440 543.200 899.560 544.320 ;
  LAYER metal3 ;
  RECT 898.440 543.200 899.560 544.320 ;
  LAYER metal2 ;
  RECT 898.440 543.200 899.560 544.320 ;
  LAYER metal1 ;
  RECT 898.440 543.200 899.560 544.320 ;
 END
END DOB28
PIN DIB27
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 885.420 543.200 886.540 544.320 ;
  LAYER metal4 ;
  RECT 885.420 543.200 886.540 544.320 ;
  LAYER metal3 ;
  RECT 885.420 543.200 886.540 544.320 ;
  LAYER metal2 ;
  RECT 885.420 543.200 886.540 544.320 ;
  LAYER metal1 ;
  RECT 885.420 543.200 886.540 544.320 ;
 END
END DIB27
PIN DOB27
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 871.780 543.200 872.900 544.320 ;
  LAYER metal4 ;
  RECT 871.780 543.200 872.900 544.320 ;
  LAYER metal3 ;
  RECT 871.780 543.200 872.900 544.320 ;
  LAYER metal2 ;
  RECT 871.780 543.200 872.900 544.320 ;
  LAYER metal1 ;
  RECT 871.780 543.200 872.900 544.320 ;
 END
END DOB27
PIN DIB26
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 858.140 543.200 859.260 544.320 ;
  LAYER metal4 ;
  RECT 858.140 543.200 859.260 544.320 ;
  LAYER metal3 ;
  RECT 858.140 543.200 859.260 544.320 ;
  LAYER metal2 ;
  RECT 858.140 543.200 859.260 544.320 ;
  LAYER metal1 ;
  RECT 858.140 543.200 859.260 544.320 ;
 END
END DIB26
PIN DOB26
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 845.120 543.200 846.240 544.320 ;
  LAYER metal4 ;
  RECT 845.120 543.200 846.240 544.320 ;
  LAYER metal3 ;
  RECT 845.120 543.200 846.240 544.320 ;
  LAYER metal2 ;
  RECT 845.120 543.200 846.240 544.320 ;
  LAYER metal1 ;
  RECT 845.120 543.200 846.240 544.320 ;
 END
END DOB26
PIN DIB25
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 831.480 543.200 832.600 544.320 ;
  LAYER metal4 ;
  RECT 831.480 543.200 832.600 544.320 ;
  LAYER metal3 ;
  RECT 831.480 543.200 832.600 544.320 ;
  LAYER metal2 ;
  RECT 831.480 543.200 832.600 544.320 ;
  LAYER metal1 ;
  RECT 831.480 543.200 832.600 544.320 ;
 END
END DIB25
PIN DOB25
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 817.840 543.200 818.960 544.320 ;
  LAYER metal4 ;
  RECT 817.840 543.200 818.960 544.320 ;
  LAYER metal3 ;
  RECT 817.840 543.200 818.960 544.320 ;
  LAYER metal2 ;
  RECT 817.840 543.200 818.960 544.320 ;
  LAYER metal1 ;
  RECT 817.840 543.200 818.960 544.320 ;
 END
END DOB25
PIN DIB24
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 804.820 543.200 805.940 544.320 ;
  LAYER metal4 ;
  RECT 804.820 543.200 805.940 544.320 ;
  LAYER metal3 ;
  RECT 804.820 543.200 805.940 544.320 ;
  LAYER metal2 ;
  RECT 804.820 543.200 805.940 544.320 ;
  LAYER metal1 ;
  RECT 804.820 543.200 805.940 544.320 ;
 END
END DIB24
PIN DOB24
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 791.180 543.200 792.300 544.320 ;
  LAYER metal4 ;
  RECT 791.180 543.200 792.300 544.320 ;
  LAYER metal3 ;
  RECT 791.180 543.200 792.300 544.320 ;
  LAYER metal2 ;
  RECT 791.180 543.200 792.300 544.320 ;
  LAYER metal1 ;
  RECT 791.180 543.200 792.300 544.320 ;
 END
END DOB24
PIN DIB23
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 777.540 543.200 778.660 544.320 ;
  LAYER metal4 ;
  RECT 777.540 543.200 778.660 544.320 ;
  LAYER metal3 ;
  RECT 777.540 543.200 778.660 544.320 ;
  LAYER metal2 ;
  RECT 777.540 543.200 778.660 544.320 ;
  LAYER metal1 ;
  RECT 777.540 543.200 778.660 544.320 ;
 END
END DIB23
PIN DOB23
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 764.520 543.200 765.640 544.320 ;
  LAYER metal4 ;
  RECT 764.520 543.200 765.640 544.320 ;
  LAYER metal3 ;
  RECT 764.520 543.200 765.640 544.320 ;
  LAYER metal2 ;
  RECT 764.520 543.200 765.640 544.320 ;
  LAYER metal1 ;
  RECT 764.520 543.200 765.640 544.320 ;
 END
END DOB23
PIN DIB22
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 750.880 543.200 752.000 544.320 ;
  LAYER metal4 ;
  RECT 750.880 543.200 752.000 544.320 ;
  LAYER metal3 ;
  RECT 750.880 543.200 752.000 544.320 ;
  LAYER metal2 ;
  RECT 750.880 543.200 752.000 544.320 ;
  LAYER metal1 ;
  RECT 750.880 543.200 752.000 544.320 ;
 END
END DIB22
PIN DOB22
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 737.240 543.200 738.360 544.320 ;
  LAYER metal4 ;
  RECT 737.240 543.200 738.360 544.320 ;
  LAYER metal3 ;
  RECT 737.240 543.200 738.360 544.320 ;
  LAYER metal2 ;
  RECT 737.240 543.200 738.360 544.320 ;
  LAYER metal1 ;
  RECT 737.240 543.200 738.360 544.320 ;
 END
END DOB22
PIN DIB21
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 724.220 543.200 725.340 544.320 ;
  LAYER metal4 ;
  RECT 724.220 543.200 725.340 544.320 ;
  LAYER metal3 ;
  RECT 724.220 543.200 725.340 544.320 ;
  LAYER metal2 ;
  RECT 724.220 543.200 725.340 544.320 ;
  LAYER metal1 ;
  RECT 724.220 543.200 725.340 544.320 ;
 END
END DIB21
PIN DOB21
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 710.580 543.200 711.700 544.320 ;
  LAYER metal4 ;
  RECT 710.580 543.200 711.700 544.320 ;
  LAYER metal3 ;
  RECT 710.580 543.200 711.700 544.320 ;
  LAYER metal2 ;
  RECT 710.580 543.200 711.700 544.320 ;
  LAYER metal1 ;
  RECT 710.580 543.200 711.700 544.320 ;
 END
END DOB21
PIN DIB20
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 696.940 543.200 698.060 544.320 ;
  LAYER metal4 ;
  RECT 696.940 543.200 698.060 544.320 ;
  LAYER metal3 ;
  RECT 696.940 543.200 698.060 544.320 ;
  LAYER metal2 ;
  RECT 696.940 543.200 698.060 544.320 ;
  LAYER metal1 ;
  RECT 696.940 543.200 698.060 544.320 ;
 END
END DIB20
PIN DOB20
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 683.920 543.200 685.040 544.320 ;
  LAYER metal4 ;
  RECT 683.920 543.200 685.040 544.320 ;
  LAYER metal3 ;
  RECT 683.920 543.200 685.040 544.320 ;
  LAYER metal2 ;
  RECT 683.920 543.200 685.040 544.320 ;
  LAYER metal1 ;
  RECT 683.920 543.200 685.040 544.320 ;
 END
END DOB20
PIN DIB19
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 670.280 543.200 671.400 544.320 ;
  LAYER metal4 ;
  RECT 670.280 543.200 671.400 544.320 ;
  LAYER metal3 ;
  RECT 670.280 543.200 671.400 544.320 ;
  LAYER metal2 ;
  RECT 670.280 543.200 671.400 544.320 ;
  LAYER metal1 ;
  RECT 670.280 543.200 671.400 544.320 ;
 END
END DIB19
PIN DOB19
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 656.640 543.200 657.760 544.320 ;
  LAYER metal4 ;
  RECT 656.640 543.200 657.760 544.320 ;
  LAYER metal3 ;
  RECT 656.640 543.200 657.760 544.320 ;
  LAYER metal2 ;
  RECT 656.640 543.200 657.760 544.320 ;
  LAYER metal1 ;
  RECT 656.640 543.200 657.760 544.320 ;
 END
END DOB19
PIN DIB18
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 643.000 543.200 644.120 544.320 ;
  LAYER metal4 ;
  RECT 643.000 543.200 644.120 544.320 ;
  LAYER metal3 ;
  RECT 643.000 543.200 644.120 544.320 ;
  LAYER metal2 ;
  RECT 643.000 543.200 644.120 544.320 ;
  LAYER metal1 ;
  RECT 643.000 543.200 644.120 544.320 ;
 END
END DIB18
PIN DOB18
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 629.980 543.200 631.100 544.320 ;
  LAYER metal4 ;
  RECT 629.980 543.200 631.100 544.320 ;
  LAYER metal3 ;
  RECT 629.980 543.200 631.100 544.320 ;
  LAYER metal2 ;
  RECT 629.980 543.200 631.100 544.320 ;
  LAYER metal1 ;
  RECT 629.980 543.200 631.100 544.320 ;
 END
END DOB18
PIN DIB17
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 616.340 543.200 617.460 544.320 ;
  LAYER metal4 ;
  RECT 616.340 543.200 617.460 544.320 ;
  LAYER metal3 ;
  RECT 616.340 543.200 617.460 544.320 ;
  LAYER metal2 ;
  RECT 616.340 543.200 617.460 544.320 ;
  LAYER metal1 ;
  RECT 616.340 543.200 617.460 544.320 ;
 END
END DIB17
PIN DOB17
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 602.700 543.200 603.820 544.320 ;
  LAYER metal4 ;
  RECT 602.700 543.200 603.820 544.320 ;
  LAYER metal3 ;
  RECT 602.700 543.200 603.820 544.320 ;
  LAYER metal2 ;
  RECT 602.700 543.200 603.820 544.320 ;
  LAYER metal1 ;
  RECT 602.700 543.200 603.820 544.320 ;
 END
END DOB17
PIN DIB16
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 589.680 543.200 590.800 544.320 ;
  LAYER metal4 ;
  RECT 589.680 543.200 590.800 544.320 ;
  LAYER metal3 ;
  RECT 589.680 543.200 590.800 544.320 ;
  LAYER metal2 ;
  RECT 589.680 543.200 590.800 544.320 ;
  LAYER metal1 ;
  RECT 589.680 543.200 590.800 544.320 ;
 END
END DIB16
PIN WEBN1
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 578.520 543.200 579.640 544.320 ;
  LAYER metal4 ;
  RECT 578.520 543.200 579.640 544.320 ;
  LAYER metal3 ;
  RECT 578.520 543.200 579.640 544.320 ;
  LAYER metal2 ;
  RECT 578.520 543.200 579.640 544.320 ;
  LAYER metal1 ;
  RECT 578.520 543.200 579.640 544.320 ;
 END
END WEBN1
PIN DOB16
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 576.040 543.200 577.160 544.320 ;
  LAYER metal4 ;
  RECT 576.040 543.200 577.160 544.320 ;
  LAYER metal3 ;
  RECT 576.040 543.200 577.160 544.320 ;
  LAYER metal2 ;
  RECT 576.040 543.200 577.160 544.320 ;
  LAYER metal1 ;
  RECT 576.040 543.200 577.160 544.320 ;
 END
END DOB16
PIN OEB
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 549.380 543.200 550.500 544.320 ;
  LAYER metal4 ;
  RECT 549.380 543.200 550.500 544.320 ;
  LAYER metal3 ;
  RECT 549.380 543.200 550.500 544.320 ;
  LAYER metal2 ;
  RECT 549.380 543.200 550.500 544.320 ;
  LAYER metal1 ;
  RECT 549.380 543.200 550.500 544.320 ;
 END
END OEB
PIN CKB
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 536.360 543.200 537.480 544.320 ;
  LAYER metal4 ;
  RECT 536.360 543.200 537.480 544.320 ;
  LAYER metal3 ;
  RECT 536.360 543.200 537.480 544.320 ;
  LAYER metal2 ;
  RECT 536.360 543.200 537.480 544.320 ;
  LAYER metal1 ;
  RECT 536.360 543.200 537.480 544.320 ;
 END
END CKB
PIN CSB
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 534.500 543.200 535.620 544.320 ;
  LAYER metal4 ;
  RECT 534.500 543.200 535.620 544.320 ;
  LAYER metal3 ;
  RECT 534.500 543.200 535.620 544.320 ;
  LAYER metal2 ;
  RECT 534.500 543.200 535.620 544.320 ;
  LAYER metal1 ;
  RECT 534.500 543.200 535.620 544.320 ;
 END
END CSB
PIN B2
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 527.680 543.200 528.800 544.320 ;
  LAYER metal4 ;
  RECT 527.680 543.200 528.800 544.320 ;
  LAYER metal3 ;
  RECT 527.680 543.200 528.800 544.320 ;
  LAYER metal2 ;
  RECT 527.680 543.200 528.800 544.320 ;
  LAYER metal1 ;
  RECT 527.680 543.200 528.800 544.320 ;
 END
END B2
PIN B1
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 522.720 543.200 523.840 544.320 ;
  LAYER metal4 ;
  RECT 522.720 543.200 523.840 544.320 ;
  LAYER metal3 ;
  RECT 522.720 543.200 523.840 544.320 ;
  LAYER metal2 ;
  RECT 522.720 543.200 523.840 544.320 ;
  LAYER metal1 ;
  RECT 522.720 543.200 523.840 544.320 ;
 END
END B1
PIN B0
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 520.240 543.200 521.360 544.320 ;
  LAYER metal4 ;
  RECT 520.240 543.200 521.360 544.320 ;
  LAYER metal3 ;
  RECT 520.240 543.200 521.360 544.320 ;
  LAYER metal2 ;
  RECT 520.240 543.200 521.360 544.320 ;
  LAYER metal1 ;
  RECT 520.240 543.200 521.360 544.320 ;
 END
END B0
PIN B5
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 511.560 543.200 512.680 544.320 ;
  LAYER metal4 ;
  RECT 511.560 543.200 512.680 544.320 ;
  LAYER metal3 ;
  RECT 511.560 543.200 512.680 544.320 ;
  LAYER metal2 ;
  RECT 511.560 543.200 512.680 544.320 ;
  LAYER metal1 ;
  RECT 511.560 543.200 512.680 544.320 ;
 END
END B5
PIN B4
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 505.980 543.200 507.100 544.320 ;
  LAYER metal4 ;
  RECT 505.980 543.200 507.100 544.320 ;
  LAYER metal3 ;
  RECT 505.980 543.200 507.100 544.320 ;
  LAYER metal2 ;
  RECT 505.980 543.200 507.100 544.320 ;
  LAYER metal1 ;
  RECT 505.980 543.200 507.100 544.320 ;
 END
END B4
PIN B3
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 500.400 543.200 501.520 544.320 ;
  LAYER metal4 ;
  RECT 500.400 543.200 501.520 544.320 ;
  LAYER metal3 ;
  RECT 500.400 543.200 501.520 544.320 ;
  LAYER metal2 ;
  RECT 500.400 543.200 501.520 544.320 ;
  LAYER metal1 ;
  RECT 500.400 543.200 501.520 544.320 ;
 END
END B3
PIN B8
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 487.380 543.200 488.500 544.320 ;
  LAYER metal4 ;
  RECT 487.380 543.200 488.500 544.320 ;
  LAYER metal3 ;
  RECT 487.380 543.200 488.500 544.320 ;
  LAYER metal2 ;
  RECT 487.380 543.200 488.500 544.320 ;
  LAYER metal1 ;
  RECT 487.380 543.200 488.500 544.320 ;
 END
END B8
PIN B7
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 481.800 543.200 482.920 544.320 ;
  LAYER metal4 ;
  RECT 481.800 543.200 482.920 544.320 ;
  LAYER metal3 ;
  RECT 481.800 543.200 482.920 544.320 ;
  LAYER metal2 ;
  RECT 481.800 543.200 482.920 544.320 ;
  LAYER metal1 ;
  RECT 481.800 543.200 482.920 544.320 ;
 END
END B7
PIN B6
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 476.220 543.200 477.340 544.320 ;
  LAYER metal4 ;
  RECT 476.220 543.200 477.340 544.320 ;
  LAYER metal3 ;
  RECT 476.220 543.200 477.340 544.320 ;
  LAYER metal2 ;
  RECT 476.220 543.200 477.340 544.320 ;
  LAYER metal1 ;
  RECT 476.220 543.200 477.340 544.320 ;
 END
END B6
PIN B9
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 451.420 543.200 452.540 544.320 ;
  LAYER metal4 ;
  RECT 451.420 543.200 452.540 544.320 ;
  LAYER metal3 ;
  RECT 451.420 543.200 452.540 544.320 ;
  LAYER metal2 ;
  RECT 451.420 543.200 452.540 544.320 ;
  LAYER metal1 ;
  RECT 451.420 543.200 452.540 544.320 ;
 END
END B9
PIN DIB15
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 429.100 543.200 430.220 544.320 ;
  LAYER metal4 ;
  RECT 429.100 543.200 430.220 544.320 ;
  LAYER metal3 ;
  RECT 429.100 543.200 430.220 544.320 ;
  LAYER metal2 ;
  RECT 429.100 543.200 430.220 544.320 ;
  LAYER metal1 ;
  RECT 429.100 543.200 430.220 544.320 ;
 END
END DIB15
PIN DOB15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 416.080 543.200 417.200 544.320 ;
  LAYER metal4 ;
  RECT 416.080 543.200 417.200 544.320 ;
  LAYER metal3 ;
  RECT 416.080 543.200 417.200 544.320 ;
  LAYER metal2 ;
  RECT 416.080 543.200 417.200 544.320 ;
  LAYER metal1 ;
  RECT 416.080 543.200 417.200 544.320 ;
 END
END DOB15
PIN DIB14
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 402.440 543.200 403.560 544.320 ;
  LAYER metal4 ;
  RECT 402.440 543.200 403.560 544.320 ;
  LAYER metal3 ;
  RECT 402.440 543.200 403.560 544.320 ;
  LAYER metal2 ;
  RECT 402.440 543.200 403.560 544.320 ;
  LAYER metal1 ;
  RECT 402.440 543.200 403.560 544.320 ;
 END
END DIB14
PIN DOB14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 388.800 543.200 389.920 544.320 ;
  LAYER metal4 ;
  RECT 388.800 543.200 389.920 544.320 ;
  LAYER metal3 ;
  RECT 388.800 543.200 389.920 544.320 ;
  LAYER metal2 ;
  RECT 388.800 543.200 389.920 544.320 ;
  LAYER metal1 ;
  RECT 388.800 543.200 389.920 544.320 ;
 END
END DOB14
PIN DIB13
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 375.780 543.200 376.900 544.320 ;
  LAYER metal4 ;
  RECT 375.780 543.200 376.900 544.320 ;
  LAYER metal3 ;
  RECT 375.780 543.200 376.900 544.320 ;
  LAYER metal2 ;
  RECT 375.780 543.200 376.900 544.320 ;
  LAYER metal1 ;
  RECT 375.780 543.200 376.900 544.320 ;
 END
END DIB13
PIN DOB13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 362.140 543.200 363.260 544.320 ;
  LAYER metal4 ;
  RECT 362.140 543.200 363.260 544.320 ;
  LAYER metal3 ;
  RECT 362.140 543.200 363.260 544.320 ;
  LAYER metal2 ;
  RECT 362.140 543.200 363.260 544.320 ;
  LAYER metal1 ;
  RECT 362.140 543.200 363.260 544.320 ;
 END
END DOB13
PIN DIB12
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 348.500 543.200 349.620 544.320 ;
  LAYER metal4 ;
  RECT 348.500 543.200 349.620 544.320 ;
  LAYER metal3 ;
  RECT 348.500 543.200 349.620 544.320 ;
  LAYER metal2 ;
  RECT 348.500 543.200 349.620 544.320 ;
  LAYER metal1 ;
  RECT 348.500 543.200 349.620 544.320 ;
 END
END DIB12
PIN DOB12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 335.480 543.200 336.600 544.320 ;
  LAYER metal4 ;
  RECT 335.480 543.200 336.600 544.320 ;
  LAYER metal3 ;
  RECT 335.480 543.200 336.600 544.320 ;
  LAYER metal2 ;
  RECT 335.480 543.200 336.600 544.320 ;
  LAYER metal1 ;
  RECT 335.480 543.200 336.600 544.320 ;
 END
END DOB12
PIN DIB11
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 321.840 543.200 322.960 544.320 ;
  LAYER metal4 ;
  RECT 321.840 543.200 322.960 544.320 ;
  LAYER metal3 ;
  RECT 321.840 543.200 322.960 544.320 ;
  LAYER metal2 ;
  RECT 321.840 543.200 322.960 544.320 ;
  LAYER metal1 ;
  RECT 321.840 543.200 322.960 544.320 ;
 END
END DIB11
PIN DOB11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 308.200 543.200 309.320 544.320 ;
  LAYER metal4 ;
  RECT 308.200 543.200 309.320 544.320 ;
  LAYER metal3 ;
  RECT 308.200 543.200 309.320 544.320 ;
  LAYER metal2 ;
  RECT 308.200 543.200 309.320 544.320 ;
  LAYER metal1 ;
  RECT 308.200 543.200 309.320 544.320 ;
 END
END DOB11
PIN DIB10
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 295.180 543.200 296.300 544.320 ;
  LAYER metal4 ;
  RECT 295.180 543.200 296.300 544.320 ;
  LAYER metal3 ;
  RECT 295.180 543.200 296.300 544.320 ;
  LAYER metal2 ;
  RECT 295.180 543.200 296.300 544.320 ;
  LAYER metal1 ;
  RECT 295.180 543.200 296.300 544.320 ;
 END
END DIB10
PIN DOB10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 281.540 543.200 282.660 544.320 ;
  LAYER metal4 ;
  RECT 281.540 543.200 282.660 544.320 ;
  LAYER metal3 ;
  RECT 281.540 543.200 282.660 544.320 ;
  LAYER metal2 ;
  RECT 281.540 543.200 282.660 544.320 ;
  LAYER metal1 ;
  RECT 281.540 543.200 282.660 544.320 ;
 END
END DOB10
PIN DIB9
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 267.900 543.200 269.020 544.320 ;
  LAYER metal4 ;
  RECT 267.900 543.200 269.020 544.320 ;
  LAYER metal3 ;
  RECT 267.900 543.200 269.020 544.320 ;
  LAYER metal2 ;
  RECT 267.900 543.200 269.020 544.320 ;
  LAYER metal1 ;
  RECT 267.900 543.200 269.020 544.320 ;
 END
END DIB9
PIN DOB9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 254.880 543.200 256.000 544.320 ;
  LAYER metal4 ;
  RECT 254.880 543.200 256.000 544.320 ;
  LAYER metal3 ;
  RECT 254.880 543.200 256.000 544.320 ;
  LAYER metal2 ;
  RECT 254.880 543.200 256.000 544.320 ;
  LAYER metal1 ;
  RECT 254.880 543.200 256.000 544.320 ;
 END
END DOB9
PIN DIB8
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 241.240 543.200 242.360 544.320 ;
  LAYER metal4 ;
  RECT 241.240 543.200 242.360 544.320 ;
  LAYER metal3 ;
  RECT 241.240 543.200 242.360 544.320 ;
  LAYER metal2 ;
  RECT 241.240 543.200 242.360 544.320 ;
  LAYER metal1 ;
  RECT 241.240 543.200 242.360 544.320 ;
 END
END DIB8
PIN DOB8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 227.600 543.200 228.720 544.320 ;
  LAYER metal4 ;
  RECT 227.600 543.200 228.720 544.320 ;
  LAYER metal3 ;
  RECT 227.600 543.200 228.720 544.320 ;
  LAYER metal2 ;
  RECT 227.600 543.200 228.720 544.320 ;
  LAYER metal1 ;
  RECT 227.600 543.200 228.720 544.320 ;
 END
END DOB8
PIN DIB7
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 214.580 543.200 215.700 544.320 ;
  LAYER metal4 ;
  RECT 214.580 543.200 215.700 544.320 ;
  LAYER metal3 ;
  RECT 214.580 543.200 215.700 544.320 ;
  LAYER metal2 ;
  RECT 214.580 543.200 215.700 544.320 ;
  LAYER metal1 ;
  RECT 214.580 543.200 215.700 544.320 ;
 END
END DIB7
PIN DOB7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 200.940 543.200 202.060 544.320 ;
  LAYER metal4 ;
  RECT 200.940 543.200 202.060 544.320 ;
  LAYER metal3 ;
  RECT 200.940 543.200 202.060 544.320 ;
  LAYER metal2 ;
  RECT 200.940 543.200 202.060 544.320 ;
  LAYER metal1 ;
  RECT 200.940 543.200 202.060 544.320 ;
 END
END DOB7
PIN DIB6
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 187.300 543.200 188.420 544.320 ;
  LAYER metal4 ;
  RECT 187.300 543.200 188.420 544.320 ;
  LAYER metal3 ;
  RECT 187.300 543.200 188.420 544.320 ;
  LAYER metal2 ;
  RECT 187.300 543.200 188.420 544.320 ;
  LAYER metal1 ;
  RECT 187.300 543.200 188.420 544.320 ;
 END
END DIB6
PIN DOB6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 174.280 543.200 175.400 544.320 ;
  LAYER metal4 ;
  RECT 174.280 543.200 175.400 544.320 ;
  LAYER metal3 ;
  RECT 174.280 543.200 175.400 544.320 ;
  LAYER metal2 ;
  RECT 174.280 543.200 175.400 544.320 ;
  LAYER metal1 ;
  RECT 174.280 543.200 175.400 544.320 ;
 END
END DOB6
PIN DIB5
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 160.640 543.200 161.760 544.320 ;
  LAYER metal4 ;
  RECT 160.640 543.200 161.760 544.320 ;
  LAYER metal3 ;
  RECT 160.640 543.200 161.760 544.320 ;
  LAYER metal2 ;
  RECT 160.640 543.200 161.760 544.320 ;
  LAYER metal1 ;
  RECT 160.640 543.200 161.760 544.320 ;
 END
END DIB5
PIN DOB5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 147.000 543.200 148.120 544.320 ;
  LAYER metal4 ;
  RECT 147.000 543.200 148.120 544.320 ;
  LAYER metal3 ;
  RECT 147.000 543.200 148.120 544.320 ;
  LAYER metal2 ;
  RECT 147.000 543.200 148.120 544.320 ;
  LAYER metal1 ;
  RECT 147.000 543.200 148.120 544.320 ;
 END
END DOB5
PIN DIB4
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 133.980 543.200 135.100 544.320 ;
  LAYER metal4 ;
  RECT 133.980 543.200 135.100 544.320 ;
  LAYER metal3 ;
  RECT 133.980 543.200 135.100 544.320 ;
  LAYER metal2 ;
  RECT 133.980 543.200 135.100 544.320 ;
  LAYER metal1 ;
  RECT 133.980 543.200 135.100 544.320 ;
 END
END DIB4
PIN DOB4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 120.340 543.200 121.460 544.320 ;
  LAYER metal4 ;
  RECT 120.340 543.200 121.460 544.320 ;
  LAYER metal3 ;
  RECT 120.340 543.200 121.460 544.320 ;
  LAYER metal2 ;
  RECT 120.340 543.200 121.460 544.320 ;
  LAYER metal1 ;
  RECT 120.340 543.200 121.460 544.320 ;
 END
END DOB4
PIN DIB3
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 106.700 543.200 107.820 544.320 ;
  LAYER metal4 ;
  RECT 106.700 543.200 107.820 544.320 ;
  LAYER metal3 ;
  RECT 106.700 543.200 107.820 544.320 ;
  LAYER metal2 ;
  RECT 106.700 543.200 107.820 544.320 ;
  LAYER metal1 ;
  RECT 106.700 543.200 107.820 544.320 ;
 END
END DIB3
PIN DOB3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 93.680 543.200 94.800 544.320 ;
  LAYER metal4 ;
  RECT 93.680 543.200 94.800 544.320 ;
  LAYER metal3 ;
  RECT 93.680 543.200 94.800 544.320 ;
  LAYER metal2 ;
  RECT 93.680 543.200 94.800 544.320 ;
  LAYER metal1 ;
  RECT 93.680 543.200 94.800 544.320 ;
 END
END DOB3
PIN DIB2
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 80.040 543.200 81.160 544.320 ;
  LAYER metal4 ;
  RECT 80.040 543.200 81.160 544.320 ;
  LAYER metal3 ;
  RECT 80.040 543.200 81.160 544.320 ;
  LAYER metal2 ;
  RECT 80.040 543.200 81.160 544.320 ;
  LAYER metal1 ;
  RECT 80.040 543.200 81.160 544.320 ;
 END
END DIB2
PIN DOB2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 66.400 543.200 67.520 544.320 ;
  LAYER metal4 ;
  RECT 66.400 543.200 67.520 544.320 ;
  LAYER metal3 ;
  RECT 66.400 543.200 67.520 544.320 ;
  LAYER metal2 ;
  RECT 66.400 543.200 67.520 544.320 ;
  LAYER metal1 ;
  RECT 66.400 543.200 67.520 544.320 ;
 END
END DOB2
PIN DIB1
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 52.760 543.200 53.880 544.320 ;
  LAYER metal4 ;
  RECT 52.760 543.200 53.880 544.320 ;
  LAYER metal3 ;
  RECT 52.760 543.200 53.880 544.320 ;
  LAYER metal2 ;
  RECT 52.760 543.200 53.880 544.320 ;
  LAYER metal1 ;
  RECT 52.760 543.200 53.880 544.320 ;
 END
END DIB1
PIN DOB1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 39.740 543.200 40.860 544.320 ;
  LAYER metal4 ;
  RECT 39.740 543.200 40.860 544.320 ;
  LAYER metal3 ;
  RECT 39.740 543.200 40.860 544.320 ;
  LAYER metal2 ;
  RECT 39.740 543.200 40.860 544.320 ;
  LAYER metal1 ;
  RECT 39.740 543.200 40.860 544.320 ;
 END
END DOB1
PIN DIB0
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 26.100 543.200 27.220 544.320 ;
  LAYER metal4 ;
  RECT 26.100 543.200 27.220 544.320 ;
  LAYER metal3 ;
  RECT 26.100 543.200 27.220 544.320 ;
  LAYER metal2 ;
  RECT 26.100 543.200 27.220 544.320 ;
  LAYER metal1 ;
  RECT 26.100 543.200 27.220 544.320 ;
 END
END DIB0
PIN WEBN0
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 14.940 543.200 16.060 544.320 ;
  LAYER metal4 ;
  RECT 14.940 543.200 16.060 544.320 ;
  LAYER metal3 ;
  RECT 14.940 543.200 16.060 544.320 ;
  LAYER metal2 ;
  RECT 14.940 543.200 16.060 544.320 ;
  LAYER metal1 ;
  RECT 14.940 543.200 16.060 544.320 ;
 END
END WEBN0
PIN DOB0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 12.460 543.200 13.580 544.320 ;
  LAYER metal4 ;
  RECT 12.460 543.200 13.580 544.320 ;
  LAYER metal3 ;
  RECT 12.460 543.200 13.580 544.320 ;
  LAYER metal2 ;
  RECT 12.460 543.200 13.580 544.320 ;
  LAYER metal1 ;
  RECT 12.460 543.200 13.580 544.320 ;
 END
END DOB0
PIN DIA47
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1422.960 0.000 1424.080 1.120 ;
  LAYER metal4 ;
  RECT 1422.960 0.000 1424.080 1.120 ;
  LAYER metal3 ;
  RECT 1422.960 0.000 1424.080 1.120 ;
  LAYER metal2 ;
  RECT 1422.960 0.000 1424.080 1.120 ;
  LAYER metal1 ;
  RECT 1422.960 0.000 1424.080 1.120 ;
 END
END DIA47
PIN DOA47
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1409.320 0.000 1410.440 1.120 ;
  LAYER metal4 ;
  RECT 1409.320 0.000 1410.440 1.120 ;
  LAYER metal3 ;
  RECT 1409.320 0.000 1410.440 1.120 ;
  LAYER metal2 ;
  RECT 1409.320 0.000 1410.440 1.120 ;
  LAYER metal1 ;
  RECT 1409.320 0.000 1410.440 1.120 ;
 END
END DOA47
PIN DIA46
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1395.680 0.000 1396.800 1.120 ;
  LAYER metal4 ;
  RECT 1395.680 0.000 1396.800 1.120 ;
  LAYER metal3 ;
  RECT 1395.680 0.000 1396.800 1.120 ;
  LAYER metal2 ;
  RECT 1395.680 0.000 1396.800 1.120 ;
  LAYER metal1 ;
  RECT 1395.680 0.000 1396.800 1.120 ;
 END
END DIA46
PIN DOA46
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1382.660 0.000 1383.780 1.120 ;
  LAYER metal4 ;
  RECT 1382.660 0.000 1383.780 1.120 ;
  LAYER metal3 ;
  RECT 1382.660 0.000 1383.780 1.120 ;
  LAYER metal2 ;
  RECT 1382.660 0.000 1383.780 1.120 ;
  LAYER metal1 ;
  RECT 1382.660 0.000 1383.780 1.120 ;
 END
END DOA46
PIN DIA45
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1369.020 0.000 1370.140 1.120 ;
  LAYER metal4 ;
  RECT 1369.020 0.000 1370.140 1.120 ;
  LAYER metal3 ;
  RECT 1369.020 0.000 1370.140 1.120 ;
  LAYER metal2 ;
  RECT 1369.020 0.000 1370.140 1.120 ;
  LAYER metal1 ;
  RECT 1369.020 0.000 1370.140 1.120 ;
 END
END DIA45
PIN DOA45
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1355.380 0.000 1356.500 1.120 ;
  LAYER metal4 ;
  RECT 1355.380 0.000 1356.500 1.120 ;
  LAYER metal3 ;
  RECT 1355.380 0.000 1356.500 1.120 ;
  LAYER metal2 ;
  RECT 1355.380 0.000 1356.500 1.120 ;
  LAYER metal1 ;
  RECT 1355.380 0.000 1356.500 1.120 ;
 END
END DOA45
PIN DIA44
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1342.360 0.000 1343.480 1.120 ;
  LAYER metal4 ;
  RECT 1342.360 0.000 1343.480 1.120 ;
  LAYER metal3 ;
  RECT 1342.360 0.000 1343.480 1.120 ;
  LAYER metal2 ;
  RECT 1342.360 0.000 1343.480 1.120 ;
  LAYER metal1 ;
  RECT 1342.360 0.000 1343.480 1.120 ;
 END
END DIA44
PIN DOA44
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1328.720 0.000 1329.840 1.120 ;
  LAYER metal4 ;
  RECT 1328.720 0.000 1329.840 1.120 ;
  LAYER metal3 ;
  RECT 1328.720 0.000 1329.840 1.120 ;
  LAYER metal2 ;
  RECT 1328.720 0.000 1329.840 1.120 ;
  LAYER metal1 ;
  RECT 1328.720 0.000 1329.840 1.120 ;
 END
END DOA44
PIN DIA43
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1315.080 0.000 1316.200 1.120 ;
  LAYER metal4 ;
  RECT 1315.080 0.000 1316.200 1.120 ;
  LAYER metal3 ;
  RECT 1315.080 0.000 1316.200 1.120 ;
  LAYER metal2 ;
  RECT 1315.080 0.000 1316.200 1.120 ;
  LAYER metal1 ;
  RECT 1315.080 0.000 1316.200 1.120 ;
 END
END DIA43
PIN DOA43
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1302.060 0.000 1303.180 1.120 ;
  LAYER metal4 ;
  RECT 1302.060 0.000 1303.180 1.120 ;
  LAYER metal3 ;
  RECT 1302.060 0.000 1303.180 1.120 ;
  LAYER metal2 ;
  RECT 1302.060 0.000 1303.180 1.120 ;
  LAYER metal1 ;
  RECT 1302.060 0.000 1303.180 1.120 ;
 END
END DOA43
PIN DIA42
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1288.420 0.000 1289.540 1.120 ;
  LAYER metal4 ;
  RECT 1288.420 0.000 1289.540 1.120 ;
  LAYER metal3 ;
  RECT 1288.420 0.000 1289.540 1.120 ;
  LAYER metal2 ;
  RECT 1288.420 0.000 1289.540 1.120 ;
  LAYER metal1 ;
  RECT 1288.420 0.000 1289.540 1.120 ;
 END
END DIA42
PIN DOA42
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1274.780 0.000 1275.900 1.120 ;
  LAYER metal4 ;
  RECT 1274.780 0.000 1275.900 1.120 ;
  LAYER metal3 ;
  RECT 1274.780 0.000 1275.900 1.120 ;
  LAYER metal2 ;
  RECT 1274.780 0.000 1275.900 1.120 ;
  LAYER metal1 ;
  RECT 1274.780 0.000 1275.900 1.120 ;
 END
END DOA42
PIN DIA41
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1261.760 0.000 1262.880 1.120 ;
  LAYER metal4 ;
  RECT 1261.760 0.000 1262.880 1.120 ;
  LAYER metal3 ;
  RECT 1261.760 0.000 1262.880 1.120 ;
  LAYER metal2 ;
  RECT 1261.760 0.000 1262.880 1.120 ;
  LAYER metal1 ;
  RECT 1261.760 0.000 1262.880 1.120 ;
 END
END DIA41
PIN DOA41
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1248.120 0.000 1249.240 1.120 ;
  LAYER metal4 ;
  RECT 1248.120 0.000 1249.240 1.120 ;
  LAYER metal3 ;
  RECT 1248.120 0.000 1249.240 1.120 ;
  LAYER metal2 ;
  RECT 1248.120 0.000 1249.240 1.120 ;
  LAYER metal1 ;
  RECT 1248.120 0.000 1249.240 1.120 ;
 END
END DOA41
PIN DIA40
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1234.480 0.000 1235.600 1.120 ;
  LAYER metal4 ;
  RECT 1234.480 0.000 1235.600 1.120 ;
  LAYER metal3 ;
  RECT 1234.480 0.000 1235.600 1.120 ;
  LAYER metal2 ;
  RECT 1234.480 0.000 1235.600 1.120 ;
  LAYER metal1 ;
  RECT 1234.480 0.000 1235.600 1.120 ;
 END
END DIA40
PIN DOA40
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1221.460 0.000 1222.580 1.120 ;
  LAYER metal4 ;
  RECT 1221.460 0.000 1222.580 1.120 ;
  LAYER metal3 ;
  RECT 1221.460 0.000 1222.580 1.120 ;
  LAYER metal2 ;
  RECT 1221.460 0.000 1222.580 1.120 ;
  LAYER metal1 ;
  RECT 1221.460 0.000 1222.580 1.120 ;
 END
END DOA40
PIN DIA39
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1207.820 0.000 1208.940 1.120 ;
  LAYER metal4 ;
  RECT 1207.820 0.000 1208.940 1.120 ;
  LAYER metal3 ;
  RECT 1207.820 0.000 1208.940 1.120 ;
  LAYER metal2 ;
  RECT 1207.820 0.000 1208.940 1.120 ;
  LAYER metal1 ;
  RECT 1207.820 0.000 1208.940 1.120 ;
 END
END DIA39
PIN DOA39
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1194.180 0.000 1195.300 1.120 ;
  LAYER metal4 ;
  RECT 1194.180 0.000 1195.300 1.120 ;
  LAYER metal3 ;
  RECT 1194.180 0.000 1195.300 1.120 ;
  LAYER metal2 ;
  RECT 1194.180 0.000 1195.300 1.120 ;
  LAYER metal1 ;
  RECT 1194.180 0.000 1195.300 1.120 ;
 END
END DOA39
PIN DIA38
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1181.160 0.000 1182.280 1.120 ;
  LAYER metal4 ;
  RECT 1181.160 0.000 1182.280 1.120 ;
  LAYER metal3 ;
  RECT 1181.160 0.000 1182.280 1.120 ;
  LAYER metal2 ;
  RECT 1181.160 0.000 1182.280 1.120 ;
  LAYER metal1 ;
  RECT 1181.160 0.000 1182.280 1.120 ;
 END
END DIA38
PIN DOA38
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1167.520 0.000 1168.640 1.120 ;
  LAYER metal4 ;
  RECT 1167.520 0.000 1168.640 1.120 ;
  LAYER metal3 ;
  RECT 1167.520 0.000 1168.640 1.120 ;
  LAYER metal2 ;
  RECT 1167.520 0.000 1168.640 1.120 ;
  LAYER metal1 ;
  RECT 1167.520 0.000 1168.640 1.120 ;
 END
END DOA38
PIN DIA37
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1153.880 0.000 1155.000 1.120 ;
  LAYER metal4 ;
  RECT 1153.880 0.000 1155.000 1.120 ;
  LAYER metal3 ;
  RECT 1153.880 0.000 1155.000 1.120 ;
  LAYER metal2 ;
  RECT 1153.880 0.000 1155.000 1.120 ;
  LAYER metal1 ;
  RECT 1153.880 0.000 1155.000 1.120 ;
 END
END DIA37
PIN DOA37
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1140.860 0.000 1141.980 1.120 ;
  LAYER metal4 ;
  RECT 1140.860 0.000 1141.980 1.120 ;
  LAYER metal3 ;
  RECT 1140.860 0.000 1141.980 1.120 ;
  LAYER metal2 ;
  RECT 1140.860 0.000 1141.980 1.120 ;
  LAYER metal1 ;
  RECT 1140.860 0.000 1141.980 1.120 ;
 END
END DOA37
PIN DIA36
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1127.220 0.000 1128.340 1.120 ;
  LAYER metal4 ;
  RECT 1127.220 0.000 1128.340 1.120 ;
  LAYER metal3 ;
  RECT 1127.220 0.000 1128.340 1.120 ;
  LAYER metal2 ;
  RECT 1127.220 0.000 1128.340 1.120 ;
  LAYER metal1 ;
  RECT 1127.220 0.000 1128.340 1.120 ;
 END
END DIA36
PIN DOA36
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1113.580 0.000 1114.700 1.120 ;
  LAYER metal4 ;
  RECT 1113.580 0.000 1114.700 1.120 ;
  LAYER metal3 ;
  RECT 1113.580 0.000 1114.700 1.120 ;
  LAYER metal2 ;
  RECT 1113.580 0.000 1114.700 1.120 ;
  LAYER metal1 ;
  RECT 1113.580 0.000 1114.700 1.120 ;
 END
END DOA36
PIN DIA35
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1100.560 0.000 1101.680 1.120 ;
  LAYER metal4 ;
  RECT 1100.560 0.000 1101.680 1.120 ;
  LAYER metal3 ;
  RECT 1100.560 0.000 1101.680 1.120 ;
  LAYER metal2 ;
  RECT 1100.560 0.000 1101.680 1.120 ;
  LAYER metal1 ;
  RECT 1100.560 0.000 1101.680 1.120 ;
 END
END DIA35
PIN DOA35
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1086.920 0.000 1088.040 1.120 ;
  LAYER metal4 ;
  RECT 1086.920 0.000 1088.040 1.120 ;
  LAYER metal3 ;
  RECT 1086.920 0.000 1088.040 1.120 ;
  LAYER metal2 ;
  RECT 1086.920 0.000 1088.040 1.120 ;
  LAYER metal1 ;
  RECT 1086.920 0.000 1088.040 1.120 ;
 END
END DOA35
PIN DIA34
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1073.280 0.000 1074.400 1.120 ;
  LAYER metal4 ;
  RECT 1073.280 0.000 1074.400 1.120 ;
  LAYER metal3 ;
  RECT 1073.280 0.000 1074.400 1.120 ;
  LAYER metal2 ;
  RECT 1073.280 0.000 1074.400 1.120 ;
  LAYER metal1 ;
  RECT 1073.280 0.000 1074.400 1.120 ;
 END
END DIA34
PIN DOA34
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1059.640 0.000 1060.760 1.120 ;
  LAYER metal4 ;
  RECT 1059.640 0.000 1060.760 1.120 ;
  LAYER metal3 ;
  RECT 1059.640 0.000 1060.760 1.120 ;
  LAYER metal2 ;
  RECT 1059.640 0.000 1060.760 1.120 ;
  LAYER metal1 ;
  RECT 1059.640 0.000 1060.760 1.120 ;
 END
END DOA34
PIN DIA33
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1046.620 0.000 1047.740 1.120 ;
  LAYER metal4 ;
  RECT 1046.620 0.000 1047.740 1.120 ;
  LAYER metal3 ;
  RECT 1046.620 0.000 1047.740 1.120 ;
  LAYER metal2 ;
  RECT 1046.620 0.000 1047.740 1.120 ;
  LAYER metal1 ;
  RECT 1046.620 0.000 1047.740 1.120 ;
 END
END DIA33
PIN DOA33
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1032.980 0.000 1034.100 1.120 ;
  LAYER metal4 ;
  RECT 1032.980 0.000 1034.100 1.120 ;
  LAYER metal3 ;
  RECT 1032.980 0.000 1034.100 1.120 ;
  LAYER metal2 ;
  RECT 1032.980 0.000 1034.100 1.120 ;
  LAYER metal1 ;
  RECT 1032.980 0.000 1034.100 1.120 ;
 END
END DOA33
PIN DIA32
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1019.340 0.000 1020.460 1.120 ;
  LAYER metal4 ;
  RECT 1019.340 0.000 1020.460 1.120 ;
  LAYER metal3 ;
  RECT 1019.340 0.000 1020.460 1.120 ;
  LAYER metal2 ;
  RECT 1019.340 0.000 1020.460 1.120 ;
  LAYER metal1 ;
  RECT 1019.340 0.000 1020.460 1.120 ;
 END
END DIA32
PIN WEAN2
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1008.180 0.000 1009.300 1.120 ;
  LAYER metal4 ;
  RECT 1008.180 0.000 1009.300 1.120 ;
  LAYER metal3 ;
  RECT 1008.180 0.000 1009.300 1.120 ;
  LAYER metal2 ;
  RECT 1008.180 0.000 1009.300 1.120 ;
  LAYER metal1 ;
  RECT 1008.180 0.000 1009.300 1.120 ;
 END
END WEAN2
PIN DOA32
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1006.320 0.000 1007.440 1.120 ;
  LAYER metal4 ;
  RECT 1006.320 0.000 1007.440 1.120 ;
  LAYER metal3 ;
  RECT 1006.320 0.000 1007.440 1.120 ;
  LAYER metal2 ;
  RECT 1006.320 0.000 1007.440 1.120 ;
  LAYER metal1 ;
  RECT 1006.320 0.000 1007.440 1.120 ;
 END
END DOA32
PIN DIA31
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 992.680 0.000 993.800 1.120 ;
  LAYER metal4 ;
  RECT 992.680 0.000 993.800 1.120 ;
  LAYER metal3 ;
  RECT 992.680 0.000 993.800 1.120 ;
  LAYER metal2 ;
  RECT 992.680 0.000 993.800 1.120 ;
  LAYER metal1 ;
  RECT 992.680 0.000 993.800 1.120 ;
 END
END DIA31
PIN DOA31
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 979.040 0.000 980.160 1.120 ;
  LAYER metal4 ;
  RECT 979.040 0.000 980.160 1.120 ;
  LAYER metal3 ;
  RECT 979.040 0.000 980.160 1.120 ;
  LAYER metal2 ;
  RECT 979.040 0.000 980.160 1.120 ;
  LAYER metal1 ;
  RECT 979.040 0.000 980.160 1.120 ;
 END
END DOA31
PIN DIA30
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 966.020 0.000 967.140 1.120 ;
  LAYER metal4 ;
  RECT 966.020 0.000 967.140 1.120 ;
  LAYER metal3 ;
  RECT 966.020 0.000 967.140 1.120 ;
  LAYER metal2 ;
  RECT 966.020 0.000 967.140 1.120 ;
  LAYER metal1 ;
  RECT 966.020 0.000 967.140 1.120 ;
 END
END DIA30
PIN DOA30
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 952.380 0.000 953.500 1.120 ;
  LAYER metal4 ;
  RECT 952.380 0.000 953.500 1.120 ;
  LAYER metal3 ;
  RECT 952.380 0.000 953.500 1.120 ;
  LAYER metal2 ;
  RECT 952.380 0.000 953.500 1.120 ;
  LAYER metal1 ;
  RECT 952.380 0.000 953.500 1.120 ;
 END
END DOA30
PIN DIA29
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 938.740 0.000 939.860 1.120 ;
  LAYER metal4 ;
  RECT 938.740 0.000 939.860 1.120 ;
  LAYER metal3 ;
  RECT 938.740 0.000 939.860 1.120 ;
  LAYER metal2 ;
  RECT 938.740 0.000 939.860 1.120 ;
  LAYER metal1 ;
  RECT 938.740 0.000 939.860 1.120 ;
 END
END DIA29
PIN DOA29
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 925.720 0.000 926.840 1.120 ;
  LAYER metal4 ;
  RECT 925.720 0.000 926.840 1.120 ;
  LAYER metal3 ;
  RECT 925.720 0.000 926.840 1.120 ;
  LAYER metal2 ;
  RECT 925.720 0.000 926.840 1.120 ;
  LAYER metal1 ;
  RECT 925.720 0.000 926.840 1.120 ;
 END
END DOA29
PIN DIA28
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 912.080 0.000 913.200 1.120 ;
  LAYER metal4 ;
  RECT 912.080 0.000 913.200 1.120 ;
  LAYER metal3 ;
  RECT 912.080 0.000 913.200 1.120 ;
  LAYER metal2 ;
  RECT 912.080 0.000 913.200 1.120 ;
  LAYER metal1 ;
  RECT 912.080 0.000 913.200 1.120 ;
 END
END DIA28
PIN DOA28
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 898.440 0.000 899.560 1.120 ;
  LAYER metal4 ;
  RECT 898.440 0.000 899.560 1.120 ;
  LAYER metal3 ;
  RECT 898.440 0.000 899.560 1.120 ;
  LAYER metal2 ;
  RECT 898.440 0.000 899.560 1.120 ;
  LAYER metal1 ;
  RECT 898.440 0.000 899.560 1.120 ;
 END
END DOA28
PIN DIA27
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 885.420 0.000 886.540 1.120 ;
  LAYER metal4 ;
  RECT 885.420 0.000 886.540 1.120 ;
  LAYER metal3 ;
  RECT 885.420 0.000 886.540 1.120 ;
  LAYER metal2 ;
  RECT 885.420 0.000 886.540 1.120 ;
  LAYER metal1 ;
  RECT 885.420 0.000 886.540 1.120 ;
 END
END DIA27
PIN DOA27
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 871.780 0.000 872.900 1.120 ;
  LAYER metal4 ;
  RECT 871.780 0.000 872.900 1.120 ;
  LAYER metal3 ;
  RECT 871.780 0.000 872.900 1.120 ;
  LAYER metal2 ;
  RECT 871.780 0.000 872.900 1.120 ;
  LAYER metal1 ;
  RECT 871.780 0.000 872.900 1.120 ;
 END
END DOA27
PIN DIA26
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 858.140 0.000 859.260 1.120 ;
  LAYER metal4 ;
  RECT 858.140 0.000 859.260 1.120 ;
  LAYER metal3 ;
  RECT 858.140 0.000 859.260 1.120 ;
  LAYER metal2 ;
  RECT 858.140 0.000 859.260 1.120 ;
  LAYER metal1 ;
  RECT 858.140 0.000 859.260 1.120 ;
 END
END DIA26
PIN DOA26
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 845.120 0.000 846.240 1.120 ;
  LAYER metal4 ;
  RECT 845.120 0.000 846.240 1.120 ;
  LAYER metal3 ;
  RECT 845.120 0.000 846.240 1.120 ;
  LAYER metal2 ;
  RECT 845.120 0.000 846.240 1.120 ;
  LAYER metal1 ;
  RECT 845.120 0.000 846.240 1.120 ;
 END
END DOA26
PIN DIA25
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 831.480 0.000 832.600 1.120 ;
  LAYER metal4 ;
  RECT 831.480 0.000 832.600 1.120 ;
  LAYER metal3 ;
  RECT 831.480 0.000 832.600 1.120 ;
  LAYER metal2 ;
  RECT 831.480 0.000 832.600 1.120 ;
  LAYER metal1 ;
  RECT 831.480 0.000 832.600 1.120 ;
 END
END DIA25
PIN DOA25
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 817.840 0.000 818.960 1.120 ;
  LAYER metal4 ;
  RECT 817.840 0.000 818.960 1.120 ;
  LAYER metal3 ;
  RECT 817.840 0.000 818.960 1.120 ;
  LAYER metal2 ;
  RECT 817.840 0.000 818.960 1.120 ;
  LAYER metal1 ;
  RECT 817.840 0.000 818.960 1.120 ;
 END
END DOA25
PIN DIA24
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 804.820 0.000 805.940 1.120 ;
  LAYER metal4 ;
  RECT 804.820 0.000 805.940 1.120 ;
  LAYER metal3 ;
  RECT 804.820 0.000 805.940 1.120 ;
  LAYER metal2 ;
  RECT 804.820 0.000 805.940 1.120 ;
  LAYER metal1 ;
  RECT 804.820 0.000 805.940 1.120 ;
 END
END DIA24
PIN DOA24
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 791.180 0.000 792.300 1.120 ;
  LAYER metal4 ;
  RECT 791.180 0.000 792.300 1.120 ;
  LAYER metal3 ;
  RECT 791.180 0.000 792.300 1.120 ;
  LAYER metal2 ;
  RECT 791.180 0.000 792.300 1.120 ;
  LAYER metal1 ;
  RECT 791.180 0.000 792.300 1.120 ;
 END
END DOA24
PIN DIA23
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 777.540 0.000 778.660 1.120 ;
  LAYER metal4 ;
  RECT 777.540 0.000 778.660 1.120 ;
  LAYER metal3 ;
  RECT 777.540 0.000 778.660 1.120 ;
  LAYER metal2 ;
  RECT 777.540 0.000 778.660 1.120 ;
  LAYER metal1 ;
  RECT 777.540 0.000 778.660 1.120 ;
 END
END DIA23
PIN DOA23
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 764.520 0.000 765.640 1.120 ;
  LAYER metal4 ;
  RECT 764.520 0.000 765.640 1.120 ;
  LAYER metal3 ;
  RECT 764.520 0.000 765.640 1.120 ;
  LAYER metal2 ;
  RECT 764.520 0.000 765.640 1.120 ;
  LAYER metal1 ;
  RECT 764.520 0.000 765.640 1.120 ;
 END
END DOA23
PIN DIA22
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 750.880 0.000 752.000 1.120 ;
  LAYER metal4 ;
  RECT 750.880 0.000 752.000 1.120 ;
  LAYER metal3 ;
  RECT 750.880 0.000 752.000 1.120 ;
  LAYER metal2 ;
  RECT 750.880 0.000 752.000 1.120 ;
  LAYER metal1 ;
  RECT 750.880 0.000 752.000 1.120 ;
 END
END DIA22
PIN DOA22
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 737.240 0.000 738.360 1.120 ;
  LAYER metal4 ;
  RECT 737.240 0.000 738.360 1.120 ;
  LAYER metal3 ;
  RECT 737.240 0.000 738.360 1.120 ;
  LAYER metal2 ;
  RECT 737.240 0.000 738.360 1.120 ;
  LAYER metal1 ;
  RECT 737.240 0.000 738.360 1.120 ;
 END
END DOA22
PIN DIA21
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 724.220 0.000 725.340 1.120 ;
  LAYER metal4 ;
  RECT 724.220 0.000 725.340 1.120 ;
  LAYER metal3 ;
  RECT 724.220 0.000 725.340 1.120 ;
  LAYER metal2 ;
  RECT 724.220 0.000 725.340 1.120 ;
  LAYER metal1 ;
  RECT 724.220 0.000 725.340 1.120 ;
 END
END DIA21
PIN DOA21
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 710.580 0.000 711.700 1.120 ;
  LAYER metal4 ;
  RECT 710.580 0.000 711.700 1.120 ;
  LAYER metal3 ;
  RECT 710.580 0.000 711.700 1.120 ;
  LAYER metal2 ;
  RECT 710.580 0.000 711.700 1.120 ;
  LAYER metal1 ;
  RECT 710.580 0.000 711.700 1.120 ;
 END
END DOA21
PIN DIA20
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 696.940 0.000 698.060 1.120 ;
  LAYER metal4 ;
  RECT 696.940 0.000 698.060 1.120 ;
  LAYER metal3 ;
  RECT 696.940 0.000 698.060 1.120 ;
  LAYER metal2 ;
  RECT 696.940 0.000 698.060 1.120 ;
  LAYER metal1 ;
  RECT 696.940 0.000 698.060 1.120 ;
 END
END DIA20
PIN DOA20
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 683.920 0.000 685.040 1.120 ;
  LAYER metal4 ;
  RECT 683.920 0.000 685.040 1.120 ;
  LAYER metal3 ;
  RECT 683.920 0.000 685.040 1.120 ;
  LAYER metal2 ;
  RECT 683.920 0.000 685.040 1.120 ;
  LAYER metal1 ;
  RECT 683.920 0.000 685.040 1.120 ;
 END
END DOA20
PIN DIA19
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 670.280 0.000 671.400 1.120 ;
  LAYER metal4 ;
  RECT 670.280 0.000 671.400 1.120 ;
  LAYER metal3 ;
  RECT 670.280 0.000 671.400 1.120 ;
  LAYER metal2 ;
  RECT 670.280 0.000 671.400 1.120 ;
  LAYER metal1 ;
  RECT 670.280 0.000 671.400 1.120 ;
 END
END DIA19
PIN DOA19
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 656.640 0.000 657.760 1.120 ;
  LAYER metal4 ;
  RECT 656.640 0.000 657.760 1.120 ;
  LAYER metal3 ;
  RECT 656.640 0.000 657.760 1.120 ;
  LAYER metal2 ;
  RECT 656.640 0.000 657.760 1.120 ;
  LAYER metal1 ;
  RECT 656.640 0.000 657.760 1.120 ;
 END
END DOA19
PIN DIA18
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 643.000 0.000 644.120 1.120 ;
  LAYER metal4 ;
  RECT 643.000 0.000 644.120 1.120 ;
  LAYER metal3 ;
  RECT 643.000 0.000 644.120 1.120 ;
  LAYER metal2 ;
  RECT 643.000 0.000 644.120 1.120 ;
  LAYER metal1 ;
  RECT 643.000 0.000 644.120 1.120 ;
 END
END DIA18
PIN DOA18
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 629.980 0.000 631.100 1.120 ;
  LAYER metal4 ;
  RECT 629.980 0.000 631.100 1.120 ;
  LAYER metal3 ;
  RECT 629.980 0.000 631.100 1.120 ;
  LAYER metal2 ;
  RECT 629.980 0.000 631.100 1.120 ;
  LAYER metal1 ;
  RECT 629.980 0.000 631.100 1.120 ;
 END
END DOA18
PIN DIA17
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 616.340 0.000 617.460 1.120 ;
  LAYER metal4 ;
  RECT 616.340 0.000 617.460 1.120 ;
  LAYER metal3 ;
  RECT 616.340 0.000 617.460 1.120 ;
  LAYER metal2 ;
  RECT 616.340 0.000 617.460 1.120 ;
  LAYER metal1 ;
  RECT 616.340 0.000 617.460 1.120 ;
 END
END DIA17
PIN DOA17
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 602.700 0.000 603.820 1.120 ;
  LAYER metal4 ;
  RECT 602.700 0.000 603.820 1.120 ;
  LAYER metal3 ;
  RECT 602.700 0.000 603.820 1.120 ;
  LAYER metal2 ;
  RECT 602.700 0.000 603.820 1.120 ;
  LAYER metal1 ;
  RECT 602.700 0.000 603.820 1.120 ;
 END
END DOA17
PIN DIA16
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 589.680 0.000 590.800 1.120 ;
  LAYER metal4 ;
  RECT 589.680 0.000 590.800 1.120 ;
  LAYER metal3 ;
  RECT 589.680 0.000 590.800 1.120 ;
  LAYER metal2 ;
  RECT 589.680 0.000 590.800 1.120 ;
  LAYER metal1 ;
  RECT 589.680 0.000 590.800 1.120 ;
 END
END DIA16
PIN WEAN1
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 578.520 0.000 579.640 1.120 ;
  LAYER metal4 ;
  RECT 578.520 0.000 579.640 1.120 ;
  LAYER metal3 ;
  RECT 578.520 0.000 579.640 1.120 ;
  LAYER metal2 ;
  RECT 578.520 0.000 579.640 1.120 ;
  LAYER metal1 ;
  RECT 578.520 0.000 579.640 1.120 ;
 END
END WEAN1
PIN DOA16
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 576.040 0.000 577.160 1.120 ;
  LAYER metal4 ;
  RECT 576.040 0.000 577.160 1.120 ;
  LAYER metal3 ;
  RECT 576.040 0.000 577.160 1.120 ;
  LAYER metal2 ;
  RECT 576.040 0.000 577.160 1.120 ;
  LAYER metal1 ;
  RECT 576.040 0.000 577.160 1.120 ;
 END
END DOA16
PIN OEA
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 549.380 0.000 550.500 1.120 ;
  LAYER metal4 ;
  RECT 549.380 0.000 550.500 1.120 ;
  LAYER metal3 ;
  RECT 549.380 0.000 550.500 1.120 ;
  LAYER metal2 ;
  RECT 549.380 0.000 550.500 1.120 ;
  LAYER metal1 ;
  RECT 549.380 0.000 550.500 1.120 ;
 END
END OEA
PIN CKA
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 536.360 0.000 537.480 1.120 ;
  LAYER metal4 ;
  RECT 536.360 0.000 537.480 1.120 ;
  LAYER metal3 ;
  RECT 536.360 0.000 537.480 1.120 ;
  LAYER metal2 ;
  RECT 536.360 0.000 537.480 1.120 ;
  LAYER metal1 ;
  RECT 536.360 0.000 537.480 1.120 ;
 END
END CKA
PIN CSA
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 534.500 0.000 535.620 1.120 ;
  LAYER metal4 ;
  RECT 534.500 0.000 535.620 1.120 ;
  LAYER metal3 ;
  RECT 534.500 0.000 535.620 1.120 ;
  LAYER metal2 ;
  RECT 534.500 0.000 535.620 1.120 ;
  LAYER metal1 ;
  RECT 534.500 0.000 535.620 1.120 ;
 END
END CSA
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 527.680 0.000 528.800 1.120 ;
  LAYER metal4 ;
  RECT 527.680 0.000 528.800 1.120 ;
  LAYER metal3 ;
  RECT 527.680 0.000 528.800 1.120 ;
  LAYER metal2 ;
  RECT 527.680 0.000 528.800 1.120 ;
  LAYER metal1 ;
  RECT 527.680 0.000 528.800 1.120 ;
 END
END A2
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 522.720 0.000 523.840 1.120 ;
  LAYER metal4 ;
  RECT 522.720 0.000 523.840 1.120 ;
  LAYER metal3 ;
  RECT 522.720 0.000 523.840 1.120 ;
  LAYER metal2 ;
  RECT 522.720 0.000 523.840 1.120 ;
  LAYER metal1 ;
  RECT 522.720 0.000 523.840 1.120 ;
 END
END A1
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 520.240 0.000 521.360 1.120 ;
  LAYER metal4 ;
  RECT 520.240 0.000 521.360 1.120 ;
  LAYER metal3 ;
  RECT 520.240 0.000 521.360 1.120 ;
  LAYER metal2 ;
  RECT 520.240 0.000 521.360 1.120 ;
  LAYER metal1 ;
  RECT 520.240 0.000 521.360 1.120 ;
 END
END A0
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 511.560 0.000 512.680 1.120 ;
  LAYER metal4 ;
  RECT 511.560 0.000 512.680 1.120 ;
  LAYER metal3 ;
  RECT 511.560 0.000 512.680 1.120 ;
  LAYER metal2 ;
  RECT 511.560 0.000 512.680 1.120 ;
  LAYER metal1 ;
  RECT 511.560 0.000 512.680 1.120 ;
 END
END A5
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 505.980 0.000 507.100 1.120 ;
  LAYER metal4 ;
  RECT 505.980 0.000 507.100 1.120 ;
  LAYER metal3 ;
  RECT 505.980 0.000 507.100 1.120 ;
  LAYER metal2 ;
  RECT 505.980 0.000 507.100 1.120 ;
  LAYER metal1 ;
  RECT 505.980 0.000 507.100 1.120 ;
 END
END A4
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 500.400 0.000 501.520 1.120 ;
  LAYER metal4 ;
  RECT 500.400 0.000 501.520 1.120 ;
  LAYER metal3 ;
  RECT 500.400 0.000 501.520 1.120 ;
  LAYER metal2 ;
  RECT 500.400 0.000 501.520 1.120 ;
  LAYER metal1 ;
  RECT 500.400 0.000 501.520 1.120 ;
 END
END A3
PIN A8
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 487.380 0.000 488.500 1.120 ;
  LAYER metal4 ;
  RECT 487.380 0.000 488.500 1.120 ;
  LAYER metal3 ;
  RECT 487.380 0.000 488.500 1.120 ;
  LAYER metal2 ;
  RECT 487.380 0.000 488.500 1.120 ;
  LAYER metal1 ;
  RECT 487.380 0.000 488.500 1.120 ;
 END
END A8
PIN A7
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 481.800 0.000 482.920 1.120 ;
  LAYER metal4 ;
  RECT 481.800 0.000 482.920 1.120 ;
  LAYER metal3 ;
  RECT 481.800 0.000 482.920 1.120 ;
  LAYER metal2 ;
  RECT 481.800 0.000 482.920 1.120 ;
  LAYER metal1 ;
  RECT 481.800 0.000 482.920 1.120 ;
 END
END A7
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 476.220 0.000 477.340 1.120 ;
  LAYER metal4 ;
  RECT 476.220 0.000 477.340 1.120 ;
  LAYER metal3 ;
  RECT 476.220 0.000 477.340 1.120 ;
  LAYER metal2 ;
  RECT 476.220 0.000 477.340 1.120 ;
  LAYER metal1 ;
  RECT 476.220 0.000 477.340 1.120 ;
 END
END A6
PIN A9
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 451.420 0.000 452.540 1.120 ;
  LAYER metal4 ;
  RECT 451.420 0.000 452.540 1.120 ;
  LAYER metal3 ;
  RECT 451.420 0.000 452.540 1.120 ;
  LAYER metal2 ;
  RECT 451.420 0.000 452.540 1.120 ;
  LAYER metal1 ;
  RECT 451.420 0.000 452.540 1.120 ;
 END
END A9
PIN DIA15
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER metal4 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER metal3 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER metal2 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER metal1 ;
  RECT 429.100 0.000 430.220 1.120 ;
 END
END DIA15
PIN DOA15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 416.080 0.000 417.200 1.120 ;
  LAYER metal4 ;
  RECT 416.080 0.000 417.200 1.120 ;
  LAYER metal3 ;
  RECT 416.080 0.000 417.200 1.120 ;
  LAYER metal2 ;
  RECT 416.080 0.000 417.200 1.120 ;
  LAYER metal1 ;
  RECT 416.080 0.000 417.200 1.120 ;
 END
END DOA15
PIN DIA14
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER metal4 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER metal3 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER metal2 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER metal1 ;
  RECT 402.440 0.000 403.560 1.120 ;
 END
END DIA14
PIN DOA14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 388.800 0.000 389.920 1.120 ;
  LAYER metal4 ;
  RECT 388.800 0.000 389.920 1.120 ;
  LAYER metal3 ;
  RECT 388.800 0.000 389.920 1.120 ;
  LAYER metal2 ;
  RECT 388.800 0.000 389.920 1.120 ;
  LAYER metal1 ;
  RECT 388.800 0.000 389.920 1.120 ;
 END
END DOA14
PIN DIA13
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 375.780 0.000 376.900 1.120 ;
  LAYER metal4 ;
  RECT 375.780 0.000 376.900 1.120 ;
  LAYER metal3 ;
  RECT 375.780 0.000 376.900 1.120 ;
  LAYER metal2 ;
  RECT 375.780 0.000 376.900 1.120 ;
  LAYER metal1 ;
  RECT 375.780 0.000 376.900 1.120 ;
 END
END DIA13
PIN DOA13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 362.140 0.000 363.260 1.120 ;
  LAYER metal4 ;
  RECT 362.140 0.000 363.260 1.120 ;
  LAYER metal3 ;
  RECT 362.140 0.000 363.260 1.120 ;
  LAYER metal2 ;
  RECT 362.140 0.000 363.260 1.120 ;
  LAYER metal1 ;
  RECT 362.140 0.000 363.260 1.120 ;
 END
END DOA13
PIN DIA12
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER metal4 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER metal3 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER metal2 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER metal1 ;
  RECT 348.500 0.000 349.620 1.120 ;
 END
END DIA12
PIN DOA12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 335.480 0.000 336.600 1.120 ;
  LAYER metal4 ;
  RECT 335.480 0.000 336.600 1.120 ;
  LAYER metal3 ;
  RECT 335.480 0.000 336.600 1.120 ;
  LAYER metal2 ;
  RECT 335.480 0.000 336.600 1.120 ;
  LAYER metal1 ;
  RECT 335.480 0.000 336.600 1.120 ;
 END
END DOA12
PIN DIA11
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 321.840 0.000 322.960 1.120 ;
  LAYER metal4 ;
  RECT 321.840 0.000 322.960 1.120 ;
  LAYER metal3 ;
  RECT 321.840 0.000 322.960 1.120 ;
  LAYER metal2 ;
  RECT 321.840 0.000 322.960 1.120 ;
  LAYER metal1 ;
  RECT 321.840 0.000 322.960 1.120 ;
 END
END DIA11
PIN DOA11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 308.200 0.000 309.320 1.120 ;
  LAYER metal4 ;
  RECT 308.200 0.000 309.320 1.120 ;
  LAYER metal3 ;
  RECT 308.200 0.000 309.320 1.120 ;
  LAYER metal2 ;
  RECT 308.200 0.000 309.320 1.120 ;
  LAYER metal1 ;
  RECT 308.200 0.000 309.320 1.120 ;
 END
END DOA11
PIN DIA10
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 295.180 0.000 296.300 1.120 ;
  LAYER metal4 ;
  RECT 295.180 0.000 296.300 1.120 ;
  LAYER metal3 ;
  RECT 295.180 0.000 296.300 1.120 ;
  LAYER metal2 ;
  RECT 295.180 0.000 296.300 1.120 ;
  LAYER metal1 ;
  RECT 295.180 0.000 296.300 1.120 ;
 END
END DIA10
PIN DOA10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 281.540 0.000 282.660 1.120 ;
  LAYER metal4 ;
  RECT 281.540 0.000 282.660 1.120 ;
  LAYER metal3 ;
  RECT 281.540 0.000 282.660 1.120 ;
  LAYER metal2 ;
  RECT 281.540 0.000 282.660 1.120 ;
  LAYER metal1 ;
  RECT 281.540 0.000 282.660 1.120 ;
 END
END DOA10
PIN DIA9
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal4 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal3 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal2 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal1 ;
  RECT 267.900 0.000 269.020 1.120 ;
 END
END DIA9
PIN DOA9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER metal4 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER metal3 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER metal2 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER metal1 ;
  RECT 254.880 0.000 256.000 1.120 ;
 END
END DOA9
PIN DIA8
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal4 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal3 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal2 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal1 ;
  RECT 241.240 0.000 242.360 1.120 ;
 END
END DIA8
PIN DOA8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 227.600 0.000 228.720 1.120 ;
  LAYER metal4 ;
  RECT 227.600 0.000 228.720 1.120 ;
  LAYER metal3 ;
  RECT 227.600 0.000 228.720 1.120 ;
  LAYER metal2 ;
  RECT 227.600 0.000 228.720 1.120 ;
  LAYER metal1 ;
  RECT 227.600 0.000 228.720 1.120 ;
 END
END DOA8
PIN DIA7
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 214.580 0.000 215.700 1.120 ;
  LAYER metal4 ;
  RECT 214.580 0.000 215.700 1.120 ;
  LAYER metal3 ;
  RECT 214.580 0.000 215.700 1.120 ;
  LAYER metal2 ;
  RECT 214.580 0.000 215.700 1.120 ;
  LAYER metal1 ;
  RECT 214.580 0.000 215.700 1.120 ;
 END
END DIA7
PIN DOA7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 200.940 0.000 202.060 1.120 ;
  LAYER metal4 ;
  RECT 200.940 0.000 202.060 1.120 ;
  LAYER metal3 ;
  RECT 200.940 0.000 202.060 1.120 ;
  LAYER metal2 ;
  RECT 200.940 0.000 202.060 1.120 ;
  LAYER metal1 ;
  RECT 200.940 0.000 202.060 1.120 ;
 END
END DOA7
PIN DIA6
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER metal4 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER metal3 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER metal2 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER metal1 ;
  RECT 187.300 0.000 188.420 1.120 ;
 END
END DIA6
PIN DOA6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 174.280 0.000 175.400 1.120 ;
  LAYER metal4 ;
  RECT 174.280 0.000 175.400 1.120 ;
  LAYER metal3 ;
  RECT 174.280 0.000 175.400 1.120 ;
  LAYER metal2 ;
  RECT 174.280 0.000 175.400 1.120 ;
  LAYER metal1 ;
  RECT 174.280 0.000 175.400 1.120 ;
 END
END DOA6
PIN DIA5
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 160.640 0.000 161.760 1.120 ;
  LAYER metal4 ;
  RECT 160.640 0.000 161.760 1.120 ;
  LAYER metal3 ;
  RECT 160.640 0.000 161.760 1.120 ;
  LAYER metal2 ;
  RECT 160.640 0.000 161.760 1.120 ;
  LAYER metal1 ;
  RECT 160.640 0.000 161.760 1.120 ;
 END
END DIA5
PIN DOA5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 147.000 0.000 148.120 1.120 ;
  LAYER metal4 ;
  RECT 147.000 0.000 148.120 1.120 ;
  LAYER metal3 ;
  RECT 147.000 0.000 148.120 1.120 ;
  LAYER metal2 ;
  RECT 147.000 0.000 148.120 1.120 ;
  LAYER metal1 ;
  RECT 147.000 0.000 148.120 1.120 ;
 END
END DOA5
PIN DIA4
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER metal4 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER metal3 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER metal2 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER metal1 ;
  RECT 133.980 0.000 135.100 1.120 ;
 END
END DIA4
PIN DOA4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 120.340 0.000 121.460 1.120 ;
  LAYER metal4 ;
  RECT 120.340 0.000 121.460 1.120 ;
  LAYER metal3 ;
  RECT 120.340 0.000 121.460 1.120 ;
  LAYER metal2 ;
  RECT 120.340 0.000 121.460 1.120 ;
  LAYER metal1 ;
  RECT 120.340 0.000 121.460 1.120 ;
 END
END DOA4
PIN DIA3
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal4 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal3 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal2 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal1 ;
  RECT 106.700 0.000 107.820 1.120 ;
 END
END DIA3
PIN DOA3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 93.680 0.000 94.800 1.120 ;
  LAYER metal4 ;
  RECT 93.680 0.000 94.800 1.120 ;
  LAYER metal3 ;
  RECT 93.680 0.000 94.800 1.120 ;
  LAYER metal2 ;
  RECT 93.680 0.000 94.800 1.120 ;
  LAYER metal1 ;
  RECT 93.680 0.000 94.800 1.120 ;
 END
END DOA3
PIN DIA2
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 80.040 0.000 81.160 1.120 ;
  LAYER metal4 ;
  RECT 80.040 0.000 81.160 1.120 ;
  LAYER metal3 ;
  RECT 80.040 0.000 81.160 1.120 ;
  LAYER metal2 ;
  RECT 80.040 0.000 81.160 1.120 ;
  LAYER metal1 ;
  RECT 80.040 0.000 81.160 1.120 ;
 END
END DIA2
PIN DOA2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 66.400 0.000 67.520 1.120 ;
  LAYER metal4 ;
  RECT 66.400 0.000 67.520 1.120 ;
  LAYER metal3 ;
  RECT 66.400 0.000 67.520 1.120 ;
  LAYER metal2 ;
  RECT 66.400 0.000 67.520 1.120 ;
  LAYER metal1 ;
  RECT 66.400 0.000 67.520 1.120 ;
 END
END DOA2
PIN DIA1
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER metal4 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER metal3 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER metal2 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER metal1 ;
  RECT 52.760 0.000 53.880 1.120 ;
 END
END DIA1
PIN DOA1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER metal4 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER metal3 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER metal2 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER metal1 ;
  RECT 39.740 0.000 40.860 1.120 ;
 END
END DOA1
PIN DIA0
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER metal4 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER metal3 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER metal2 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER metal1 ;
  RECT 26.100 0.000 27.220 1.120 ;
 END
END DIA0
PIN WEAN0
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 14.940 0.000 16.060 1.120 ;
  LAYER metal4 ;
  RECT 14.940 0.000 16.060 1.120 ;
  LAYER metal3 ;
  RECT 14.940 0.000 16.060 1.120 ;
  LAYER metal2 ;
  RECT 14.940 0.000 16.060 1.120 ;
  LAYER metal1 ;
  RECT 14.940 0.000 16.060 1.120 ;
 END
END WEAN0
PIN DOA0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER metal4 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER metal3 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER metal2 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER metal1 ;
  RECT 12.460 0.000 13.580 1.120 ;
 END
END DOA0
OBS
  LAYER metal1 SPACING 0.280 ;
  RECT 0.000 0.140 1445.840 544.180 ;
  LAYER metal2 SPACING 0.320 ;
  RECT 0.000 0.140 1445.840 544.180 ;
  LAYER metal3 SPACING 0.320 ;
  RECT 0.000 0.140 1445.840 544.180 ;
  LAYER metal4 SPACING 0.600 ;
  RECT 0.000 0.140 1445.840 544.180 ;
  LAYER via ;
  RECT 0.000 0.140 1445.840 544.180 ;
  LAYER via2 ;
  RECT 0.000 0.140 1445.840 544.180 ;
  LAYER via3 ;
  RECT 0.000 0.140 1445.840 544.180 ;
END
END pixel_sram
END LIBRARY



