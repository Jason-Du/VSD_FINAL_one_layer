`timescale 1ns/10ps
module cnn_wrapper(

);

//bus port should wait setting state


//interrupt_output
//enable_write_interrupt signal