module cnn_top(
	clk,
	rst,
	input_data,
	predict_result
);