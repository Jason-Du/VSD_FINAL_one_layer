`timescale 1ns/10ps
module cnn_wrapper(

);

//bus port should wait setting state


//interrupt_output

//cpu clean 

//dma start